magic
tech sky130A
magscale 1 2
timestamp 1647927934
<< obsli1 >>
rect 1104 527 127420 126769
<< obsm1 >>
rect 1104 496 127420 126800
<< metal2 >>
rect 634 128302 746 129102
rect 2566 128302 2678 129102
rect 5142 128302 5254 129102
rect 7718 128302 7830 129102
rect 10294 128302 10406 129102
rect 12226 128302 12338 129102
rect 14802 128302 14914 129102
rect 17378 128302 17490 129102
rect 19310 128302 19422 129102
rect 21886 128302 21998 129102
rect 24462 128302 24574 129102
rect 26394 128302 26506 129102
rect 28970 128302 29082 129102
rect 31546 128302 31658 129102
rect 33478 128302 33590 129102
rect 36054 128302 36166 129102
rect 38630 128302 38742 129102
rect 40562 128302 40674 129102
rect 43138 128302 43250 129102
rect 45714 128302 45826 129102
rect 47646 128302 47758 129102
rect 50222 128302 50334 129102
rect 52798 128302 52910 129102
rect 54730 128302 54842 129102
rect 57306 128302 57418 129102
rect 59882 128302 59994 129102
rect 61814 128302 61926 129102
rect 64390 128302 64502 129102
rect 66966 128302 67078 129102
rect 69542 128302 69654 129102
rect 71474 128302 71586 129102
rect 74050 128302 74162 129102
rect 76626 128302 76738 129102
rect 78558 128302 78670 129102
rect 81134 128302 81246 129102
rect 83710 128302 83822 129102
rect 85642 128302 85754 129102
rect 88218 128302 88330 129102
rect 90794 128302 90906 129102
rect 92726 128302 92838 129102
rect 95302 128302 95414 129102
rect 97878 128302 97990 129102
rect 99810 128302 99922 129102
rect 102386 128302 102498 129102
rect 104962 128302 105074 129102
rect 106894 128302 107006 129102
rect 109470 128302 109582 129102
rect 112046 128302 112158 129102
rect 113978 128302 114090 129102
rect 116554 128302 116666 129102
rect 119130 128302 119242 129102
rect 121062 128302 121174 129102
rect 123638 128302 123750 129102
rect 126214 128302 126326 129102
rect 128146 128302 128258 129102
rect -10 0 102 800
rect 1922 0 2034 800
rect 4498 0 4610 800
rect 7074 0 7186 800
rect 9006 0 9118 800
rect 11582 0 11694 800
rect 14158 0 14270 800
rect 16090 0 16202 800
rect 18666 0 18778 800
rect 21242 0 21354 800
rect 23174 0 23286 800
rect 25750 0 25862 800
rect 28326 0 28438 800
rect 30258 0 30370 800
rect 32834 0 32946 800
rect 35410 0 35522 800
rect 37342 0 37454 800
rect 39918 0 40030 800
rect 42494 0 42606 800
rect 44426 0 44538 800
rect 47002 0 47114 800
rect 49578 0 49690 800
rect 51510 0 51622 800
rect 54086 0 54198 800
rect 56662 0 56774 800
rect 58594 0 58706 800
rect 61170 0 61282 800
rect 63746 0 63858 800
rect 66322 0 66434 800
rect 68254 0 68366 800
rect 70830 0 70942 800
rect 73406 0 73518 800
rect 75338 0 75450 800
rect 77914 0 78026 800
rect 80490 0 80602 800
rect 82422 0 82534 800
rect 84998 0 85110 800
rect 87574 0 87686 800
rect 89506 0 89618 800
rect 92082 0 92194 800
rect 94658 0 94770 800
rect 96590 0 96702 800
rect 99166 0 99278 800
rect 101742 0 101854 800
rect 103674 0 103786 800
rect 106250 0 106362 800
rect 108826 0 108938 800
rect 110758 0 110870 800
rect 113334 0 113446 800
rect 115910 0 116022 800
rect 117842 0 117954 800
rect 120418 0 120530 800
rect 122994 0 123106 800
rect 125570 0 125682 800
rect 127502 0 127614 800
<< obsm2 >>
rect 1398 128246 2510 128330
rect 2734 128246 5086 128330
rect 5310 128246 7662 128330
rect 7886 128246 10238 128330
rect 10462 128246 12170 128330
rect 12394 128246 14746 128330
rect 14970 128246 17322 128330
rect 17546 128246 19254 128330
rect 19478 128246 21830 128330
rect 22054 128246 24406 128330
rect 24630 128246 26338 128330
rect 26562 128246 28914 128330
rect 29138 128246 31490 128330
rect 31714 128246 33422 128330
rect 33646 128246 35998 128330
rect 36222 128246 38574 128330
rect 38798 128246 40506 128330
rect 40730 128246 43082 128330
rect 43306 128246 45658 128330
rect 45882 128246 47590 128330
rect 47814 128246 50166 128330
rect 50390 128246 52742 128330
rect 52966 128246 54674 128330
rect 54898 128246 57250 128330
rect 57474 128246 59826 128330
rect 60050 128246 61758 128330
rect 61982 128246 64334 128330
rect 64558 128246 66910 128330
rect 67134 128246 69486 128330
rect 69710 128246 71418 128330
rect 71642 128246 73994 128330
rect 74218 128246 76570 128330
rect 76794 128246 78502 128330
rect 78726 128246 81078 128330
rect 81302 128246 83654 128330
rect 83878 128246 85586 128330
rect 85810 128246 88162 128330
rect 88386 128246 90738 128330
rect 90962 128246 92670 128330
rect 92894 128246 95246 128330
rect 95470 128246 97822 128330
rect 98046 128246 99754 128330
rect 99978 128246 102330 128330
rect 102554 128246 104906 128330
rect 105130 128246 106838 128330
rect 107062 128246 109414 128330
rect 109638 128246 111990 128330
rect 112214 128246 113922 128330
rect 114146 128246 116498 128330
rect 116722 128246 119074 128330
rect 119298 128246 121006 128330
rect 121230 128246 123582 128330
rect 123806 128246 126158 128330
rect 126382 128246 126850 128330
rect 1398 856 126850 128246
rect 1398 496 1866 856
rect 2090 496 4442 856
rect 4666 496 7018 856
rect 7242 496 8950 856
rect 9174 496 11526 856
rect 11750 496 14102 856
rect 14326 496 16034 856
rect 16258 496 18610 856
rect 18834 496 21186 856
rect 21410 496 23118 856
rect 23342 496 25694 856
rect 25918 496 28270 856
rect 28494 496 30202 856
rect 30426 496 32778 856
rect 33002 496 35354 856
rect 35578 496 37286 856
rect 37510 496 39862 856
rect 40086 496 42438 856
rect 42662 496 44370 856
rect 44594 496 46946 856
rect 47170 496 49522 856
rect 49746 496 51454 856
rect 51678 496 54030 856
rect 54254 496 56606 856
rect 56830 496 58538 856
rect 58762 496 61114 856
rect 61338 496 63690 856
rect 63914 496 66266 856
rect 66490 496 68198 856
rect 68422 496 70774 856
rect 70998 496 73350 856
rect 73574 496 75282 856
rect 75506 496 77858 856
rect 78082 496 80434 856
rect 80658 496 82366 856
rect 82590 496 84942 856
rect 85166 496 87518 856
rect 87742 496 89450 856
rect 89674 496 92026 856
rect 92250 496 94602 856
rect 94826 496 96534 856
rect 96758 496 99110 856
rect 99334 496 101686 856
rect 101910 496 103618 856
rect 103842 496 106194 856
rect 106418 496 108770 856
rect 108994 496 110702 856
rect 110926 496 113278 856
rect 113502 496 115854 856
rect 116078 496 117786 856
rect 118010 496 120362 856
rect 120586 496 122938 856
rect 123162 496 125514 856
rect 125738 496 126850 856
<< metal3 >>
rect 0 127108 800 127348
rect 127790 126428 128590 126668
rect 0 124388 800 124628
rect 127790 123708 128590 123948
rect 0 122348 800 122588
rect 127790 120988 128590 121228
rect 0 119628 800 119868
rect 127790 118948 128590 119188
rect 0 116908 800 117148
rect 127790 116228 128590 116468
rect 0 114868 800 115108
rect 127790 113508 128590 113748
rect 0 112148 800 112388
rect 127790 111468 128590 111708
rect 0 109428 800 109668
rect 127790 108748 128590 108988
rect 0 107388 800 107628
rect 127790 106028 128590 106268
rect 0 104668 800 104908
rect 127790 103988 128590 104228
rect 0 101948 800 102188
rect 127790 101268 128590 101508
rect 0 99908 800 100148
rect 127790 98548 128590 98788
rect 0 97188 800 97428
rect 127790 96508 128590 96748
rect 0 94468 800 94708
rect 127790 93788 128590 94028
rect 0 92428 800 92668
rect 127790 91068 128590 91308
rect 0 89708 800 89948
rect 127790 89028 128590 89268
rect 0 86988 800 87228
rect 127790 86308 128590 86548
rect 0 84948 800 85188
rect 127790 83588 128590 83828
rect 0 82228 800 82468
rect 127790 81548 128590 81788
rect 0 79508 800 79748
rect 127790 78828 128590 79068
rect 0 77468 800 77708
rect 127790 76108 128590 76348
rect 0 74748 800 74988
rect 127790 74068 128590 74308
rect 0 72028 800 72268
rect 127790 71348 128590 71588
rect 0 69988 800 70228
rect 127790 68628 128590 68868
rect 0 67268 800 67508
rect 127790 66588 128590 66828
rect 0 64548 800 64788
rect 127790 63868 128590 64108
rect 0 61828 800 62068
rect 127790 61148 128590 61388
rect 0 59788 800 60028
rect 127790 58428 128590 58668
rect 0 57068 800 57308
rect 127790 56388 128590 56628
rect 0 54348 800 54588
rect 127790 53668 128590 53908
rect 0 52308 800 52548
rect 127790 50948 128590 51188
rect 0 49588 800 49828
rect 127790 48908 128590 49148
rect 0 46868 800 47108
rect 127790 46188 128590 46428
rect 0 44828 800 45068
rect 127790 43468 128590 43708
rect 0 42108 800 42348
rect 127790 41428 128590 41668
rect 0 39388 800 39628
rect 127790 38708 128590 38948
rect 0 37348 800 37588
rect 127790 35988 128590 36228
rect 0 34628 800 34868
rect 127790 33948 128590 34188
rect 0 31908 800 32148
rect 127790 31228 128590 31468
rect 0 29868 800 30108
rect 127790 28508 128590 28748
rect 0 27148 800 27388
rect 127790 26468 128590 26708
rect 0 24428 800 24668
rect 127790 23748 128590 23988
rect 0 22388 800 22628
rect 127790 21028 128590 21268
rect 0 19668 800 19908
rect 127790 18988 128590 19228
rect 0 16948 800 17188
rect 127790 16268 128590 16508
rect 0 14908 800 15148
rect 127790 13548 128590 13788
rect 0 12188 800 12428
rect 127790 11508 128590 11748
rect 0 9468 800 9708
rect 127790 8788 128590 9028
rect 0 7428 800 7668
rect 127790 6068 128590 6308
rect 0 4708 800 4948
rect 127790 4028 128590 4268
rect 0 1988 800 2228
rect 127790 1308 128590 1548
<< obsm3 >>
rect 800 126748 127790 126785
rect 800 126348 127710 126748
rect 800 124708 127790 126348
rect 880 124308 127790 124708
rect 800 124028 127790 124308
rect 800 123628 127710 124028
rect 800 122668 127790 123628
rect 880 122268 127790 122668
rect 800 121308 127790 122268
rect 800 120908 127710 121308
rect 800 119948 127790 120908
rect 880 119548 127790 119948
rect 800 119268 127790 119548
rect 800 118868 127710 119268
rect 800 117228 127790 118868
rect 880 116828 127790 117228
rect 800 116548 127790 116828
rect 800 116148 127710 116548
rect 800 115188 127790 116148
rect 880 114788 127790 115188
rect 800 113828 127790 114788
rect 800 113428 127710 113828
rect 800 112468 127790 113428
rect 880 112068 127790 112468
rect 800 111788 127790 112068
rect 800 111388 127710 111788
rect 800 109748 127790 111388
rect 880 109348 127790 109748
rect 800 109068 127790 109348
rect 800 108668 127710 109068
rect 800 107708 127790 108668
rect 880 107308 127790 107708
rect 800 106348 127790 107308
rect 800 105948 127710 106348
rect 800 104988 127790 105948
rect 880 104588 127790 104988
rect 800 104308 127790 104588
rect 800 103908 127710 104308
rect 800 102268 127790 103908
rect 880 101868 127790 102268
rect 800 101588 127790 101868
rect 800 101188 127710 101588
rect 800 100228 127790 101188
rect 880 99828 127790 100228
rect 800 98868 127790 99828
rect 800 98468 127710 98868
rect 800 97508 127790 98468
rect 880 97108 127790 97508
rect 800 96828 127790 97108
rect 800 96428 127710 96828
rect 800 94788 127790 96428
rect 880 94388 127790 94788
rect 800 94108 127790 94388
rect 800 93708 127710 94108
rect 800 92748 127790 93708
rect 880 92348 127790 92748
rect 800 91388 127790 92348
rect 800 90988 127710 91388
rect 800 90028 127790 90988
rect 880 89628 127790 90028
rect 800 89348 127790 89628
rect 800 88948 127710 89348
rect 800 87308 127790 88948
rect 880 86908 127790 87308
rect 800 86628 127790 86908
rect 800 86228 127710 86628
rect 800 85268 127790 86228
rect 880 84868 127790 85268
rect 800 83908 127790 84868
rect 800 83508 127710 83908
rect 800 82548 127790 83508
rect 880 82148 127790 82548
rect 800 81868 127790 82148
rect 800 81468 127710 81868
rect 800 79828 127790 81468
rect 880 79428 127790 79828
rect 800 79148 127790 79428
rect 800 78748 127710 79148
rect 800 77788 127790 78748
rect 880 77388 127790 77788
rect 800 76428 127790 77388
rect 800 76028 127710 76428
rect 800 75068 127790 76028
rect 880 74668 127790 75068
rect 800 74388 127790 74668
rect 800 73988 127710 74388
rect 800 72348 127790 73988
rect 880 71948 127790 72348
rect 800 71668 127790 71948
rect 800 71268 127710 71668
rect 800 70308 127790 71268
rect 880 69908 127790 70308
rect 800 68948 127790 69908
rect 800 68548 127710 68948
rect 800 67588 127790 68548
rect 880 67188 127790 67588
rect 800 66908 127790 67188
rect 800 66508 127710 66908
rect 800 64868 127790 66508
rect 880 64468 127790 64868
rect 800 64188 127790 64468
rect 800 63788 127710 64188
rect 800 62148 127790 63788
rect 880 61748 127790 62148
rect 800 61468 127790 61748
rect 800 61068 127710 61468
rect 800 60108 127790 61068
rect 880 59708 127790 60108
rect 800 58748 127790 59708
rect 800 58348 127710 58748
rect 800 57388 127790 58348
rect 880 56988 127790 57388
rect 800 56708 127790 56988
rect 800 56308 127710 56708
rect 800 54668 127790 56308
rect 880 54268 127790 54668
rect 800 53988 127790 54268
rect 800 53588 127710 53988
rect 800 52628 127790 53588
rect 880 52228 127790 52628
rect 800 51268 127790 52228
rect 800 50868 127710 51268
rect 800 49908 127790 50868
rect 880 49508 127790 49908
rect 800 49228 127790 49508
rect 800 48828 127710 49228
rect 800 47188 127790 48828
rect 880 46788 127790 47188
rect 800 46508 127790 46788
rect 800 46108 127710 46508
rect 800 45148 127790 46108
rect 880 44748 127790 45148
rect 800 43788 127790 44748
rect 800 43388 127710 43788
rect 800 42428 127790 43388
rect 880 42028 127790 42428
rect 800 41748 127790 42028
rect 800 41348 127710 41748
rect 800 39708 127790 41348
rect 880 39308 127790 39708
rect 800 39028 127790 39308
rect 800 38628 127710 39028
rect 800 37668 127790 38628
rect 880 37268 127790 37668
rect 800 36308 127790 37268
rect 800 35908 127710 36308
rect 800 34948 127790 35908
rect 880 34548 127790 34948
rect 800 34268 127790 34548
rect 800 33868 127710 34268
rect 800 32228 127790 33868
rect 880 31828 127790 32228
rect 800 31548 127790 31828
rect 800 31148 127710 31548
rect 800 30188 127790 31148
rect 880 29788 127790 30188
rect 800 28828 127790 29788
rect 800 28428 127710 28828
rect 800 27468 127790 28428
rect 880 27068 127790 27468
rect 800 26788 127790 27068
rect 800 26388 127710 26788
rect 800 24748 127790 26388
rect 880 24348 127790 24748
rect 800 24068 127790 24348
rect 800 23668 127710 24068
rect 800 22708 127790 23668
rect 880 22308 127790 22708
rect 800 21348 127790 22308
rect 800 20948 127710 21348
rect 800 19988 127790 20948
rect 880 19588 127790 19988
rect 800 19308 127790 19588
rect 800 18908 127710 19308
rect 800 17268 127790 18908
rect 880 16868 127790 17268
rect 800 16588 127790 16868
rect 800 16188 127710 16588
rect 800 15228 127790 16188
rect 880 14828 127790 15228
rect 800 13868 127790 14828
rect 800 13468 127710 13868
rect 800 12508 127790 13468
rect 880 12108 127790 12508
rect 800 11828 127790 12108
rect 800 11428 127710 11828
rect 800 9788 127790 11428
rect 880 9388 127790 9788
rect 800 9108 127790 9388
rect 800 8708 127710 9108
rect 800 7748 127790 8708
rect 880 7348 127790 7748
rect 800 6388 127790 7348
rect 800 5988 127710 6388
rect 800 5028 127790 5988
rect 880 4628 127790 5028
rect 800 4348 127790 4628
rect 800 3948 127710 4348
rect 800 2308 127790 3948
rect 880 1908 127790 2308
rect 800 1628 127790 1908
rect 800 1228 127710 1628
rect 800 511 127790 1228
<< metal4 >>
rect 4208 496 4528 126800
rect 19568 496 19888 126800
rect 34928 496 35248 126800
rect 50288 496 50608 126800
rect 65648 496 65968 126800
rect 81008 496 81328 126800
rect 96368 496 96688 126800
rect 111728 496 112048 126800
<< obsm4 >>
rect 34651 14451 34848 124269
rect 35328 14451 50208 124269
rect 50688 14451 65568 124269
rect 66048 14451 80928 124269
rect 81408 14451 96288 124269
rect 96768 14451 111648 124269
rect 112128 14451 112181 124269
<< labels >>
rlabel metal3 s 0 119628 800 119868 6 active
port 1 nsew signal input
rlabel metal2 s 39918 0 40030 800 6 io_in[0]
port 2 nsew signal input
rlabel metal2 s 71474 128302 71586 129102 6 io_in[10]
port 3 nsew signal input
rlabel metal2 s 634 128302 746 129102 6 io_in[11]
port 4 nsew signal input
rlabel metal3 s 127790 108748 128590 108988 6 io_in[12]
port 5 nsew signal input
rlabel metal2 s 61170 0 61282 800 6 io_in[13]
port 6 nsew signal input
rlabel metal2 s 47646 128302 47758 129102 6 io_in[14]
port 7 nsew signal input
rlabel metal3 s 127790 113508 128590 113748 6 io_in[15]
port 8 nsew signal input
rlabel metal3 s 127790 11508 128590 11748 6 io_in[16]
port 9 nsew signal input
rlabel metal2 s 26394 128302 26506 129102 6 io_in[17]
port 10 nsew signal input
rlabel metal2 s 31546 128302 31658 129102 6 io_in[18]
port 11 nsew signal input
rlabel metal2 s 110758 0 110870 800 6 io_in[19]
port 12 nsew signal input
rlabel metal3 s 0 42108 800 42348 6 io_in[1]
port 13 nsew signal input
rlabel metal3 s 0 74748 800 74988 6 io_in[20]
port 14 nsew signal input
rlabel metal3 s 0 49588 800 49828 6 io_in[21]
port 15 nsew signal input
rlabel metal3 s 127790 41428 128590 41668 6 io_in[22]
port 16 nsew signal input
rlabel metal2 s 24462 128302 24574 129102 6 io_in[23]
port 17 nsew signal input
rlabel metal2 s 17378 128302 17490 129102 6 io_in[24]
port 18 nsew signal input
rlabel metal2 s 96590 0 96702 800 6 io_in[25]
port 19 nsew signal input
rlabel metal2 s 94658 0 94770 800 6 io_in[26]
port 20 nsew signal input
rlabel metal3 s 127790 28508 128590 28748 6 io_in[27]
port 21 nsew signal input
rlabel metal2 s 84998 0 85110 800 6 io_in[28]
port 22 nsew signal input
rlabel metal2 s 128146 128302 128258 129102 6 io_in[29]
port 23 nsew signal input
rlabel metal2 s 42494 0 42606 800 6 io_in[2]
port 24 nsew signal input
rlabel metal3 s 127790 50948 128590 51188 6 io_in[30]
port 25 nsew signal input
rlabel metal3 s 0 114868 800 115108 6 io_in[31]
port 26 nsew signal input
rlabel metal2 s 80490 0 80602 800 6 io_in[32]
port 27 nsew signal input
rlabel metal3 s 0 67268 800 67508 6 io_in[33]
port 28 nsew signal input
rlabel metal2 s 97878 128302 97990 129102 6 io_in[34]
port 29 nsew signal input
rlabel metal2 s 112046 128302 112158 129102 6 io_in[35]
port 30 nsew signal input
rlabel metal3 s 127790 81548 128590 81788 6 io_in[36]
port 31 nsew signal input
rlabel metal2 s 113978 128302 114090 129102 6 io_in[37]
port 32 nsew signal input
rlabel metal2 s 74050 128302 74162 129102 6 io_in[3]
port 33 nsew signal input
rlabel metal3 s 127790 78828 128590 79068 6 io_in[4]
port 34 nsew signal input
rlabel metal3 s 127790 123708 128590 123948 6 io_in[5]
port 35 nsew signal input
rlabel metal3 s 0 79508 800 79748 6 io_in[6]
port 36 nsew signal input
rlabel metal3 s 0 54348 800 54588 6 io_in[7]
port 37 nsew signal input
rlabel metal3 s 127790 86308 128590 86548 6 io_in[8]
port 38 nsew signal input
rlabel metal2 s 21886 128302 21998 129102 6 io_in[9]
port 39 nsew signal input
rlabel metal2 s 68254 0 68366 800 6 io_oeb[0]
port 40 nsew signal output
rlabel metal3 s 0 44828 800 45068 6 io_oeb[10]
port 41 nsew signal output
rlabel metal3 s 127790 74068 128590 74308 6 io_oeb[11]
port 42 nsew signal output
rlabel metal3 s 127790 38708 128590 38948 6 io_oeb[12]
port 43 nsew signal output
rlabel metal3 s 127790 35988 128590 36228 6 io_oeb[13]
port 44 nsew signal output
rlabel metal3 s 0 12188 800 12428 6 io_oeb[14]
port 45 nsew signal output
rlabel metal2 s 36054 128302 36166 129102 6 io_oeb[15]
port 46 nsew signal output
rlabel metal3 s 127790 6068 128590 6308 6 io_oeb[16]
port 47 nsew signal output
rlabel metal2 s 35410 0 35522 800 6 io_oeb[17]
port 48 nsew signal output
rlabel metal2 s 92726 128302 92838 129102 6 io_oeb[18]
port 49 nsew signal output
rlabel metal2 s 38630 128302 38742 129102 6 io_oeb[19]
port 50 nsew signal output
rlabel metal2 s 101742 0 101854 800 6 io_oeb[1]
port 51 nsew signal output
rlabel metal3 s 127790 56388 128590 56628 6 io_oeb[20]
port 52 nsew signal output
rlabel metal2 s 5142 128302 5254 129102 6 io_oeb[21]
port 53 nsew signal output
rlabel metal2 s 14158 0 14270 800 6 io_oeb[22]
port 54 nsew signal output
rlabel metal2 s 64390 128302 64502 129102 6 io_oeb[23]
port 55 nsew signal output
rlabel metal2 s 66966 128302 67078 129102 6 io_oeb[24]
port 56 nsew signal output
rlabel metal2 s 122994 0 123106 800 6 io_oeb[25]
port 57 nsew signal output
rlabel metal3 s 127790 101268 128590 101508 6 io_oeb[26]
port 58 nsew signal output
rlabel metal2 s 76626 128302 76738 129102 6 io_oeb[27]
port 59 nsew signal output
rlabel metal2 s 108826 0 108938 800 6 io_oeb[28]
port 60 nsew signal output
rlabel metal3 s 127790 83588 128590 83828 6 io_oeb[29]
port 61 nsew signal output
rlabel metal2 s 106894 128302 107006 129102 6 io_oeb[2]
port 62 nsew signal output
rlabel metal2 s 7718 128302 7830 129102 6 io_oeb[30]
port 63 nsew signal output
rlabel metal2 s 106250 0 106362 800 6 io_oeb[31]
port 64 nsew signal output
rlabel metal3 s 0 64548 800 64788 6 io_oeb[32]
port 65 nsew signal output
rlabel metal2 s 125570 0 125682 800 6 io_oeb[33]
port 66 nsew signal output
rlabel metal2 s 28970 128302 29082 129102 6 io_oeb[34]
port 67 nsew signal output
rlabel metal3 s 0 57068 800 57308 6 io_oeb[35]
port 68 nsew signal output
rlabel metal3 s 0 29868 800 30108 6 io_oeb[36]
port 69 nsew signal output
rlabel metal3 s 0 46868 800 47108 6 io_oeb[37]
port 70 nsew signal output
rlabel metal2 s 66322 0 66434 800 6 io_oeb[3]
port 71 nsew signal output
rlabel metal3 s 127790 1308 128590 1548 6 io_oeb[4]
port 72 nsew signal output
rlabel metal3 s 0 84948 800 85188 6 io_oeb[5]
port 73 nsew signal output
rlabel metal3 s 127790 46188 128590 46428 6 io_oeb[6]
port 74 nsew signal output
rlabel metal2 s 33478 128302 33590 129102 6 io_oeb[7]
port 75 nsew signal output
rlabel metal2 s 11582 0 11694 800 6 io_oeb[8]
port 76 nsew signal output
rlabel metal2 s 28326 0 28438 800 6 io_oeb[9]
port 77 nsew signal output
rlabel metal3 s 127790 120988 128590 121228 6 io_out[0]
port 78 nsew signal output
rlabel metal3 s 127790 71348 128590 71588 6 io_out[10]
port 79 nsew signal output
rlabel metal3 s 0 7428 800 7668 6 io_out[11]
port 80 nsew signal output
rlabel metal3 s 0 19668 800 19908 6 io_out[12]
port 81 nsew signal output
rlabel metal2 s 103674 0 103786 800 6 io_out[13]
port 82 nsew signal output
rlabel metal3 s 127790 103988 128590 104228 6 io_out[14]
port 83 nsew signal output
rlabel metal3 s 0 107388 800 107628 6 io_out[15]
port 84 nsew signal output
rlabel metal3 s 127790 68628 128590 68868 6 io_out[16]
port 85 nsew signal output
rlabel metal2 s 119130 128302 119242 129102 6 io_out[17]
port 86 nsew signal output
rlabel metal2 s 120418 0 120530 800 6 io_out[18]
port 87 nsew signal output
rlabel metal3 s 0 61828 800 62068 6 io_out[19]
port 88 nsew signal output
rlabel metal2 s 85642 128302 85754 129102 6 io_out[1]
port 89 nsew signal output
rlabel metal2 s 104962 128302 105074 129102 6 io_out[20]
port 90 nsew signal output
rlabel metal3 s 0 104668 800 104908 6 io_out[21]
port 91 nsew signal output
rlabel metal2 s 82422 0 82534 800 6 io_out[22]
port 92 nsew signal output
rlabel metal3 s 127790 58428 128590 58668 6 io_out[23]
port 93 nsew signal output
rlabel metal2 s 70830 0 70942 800 6 io_out[24]
port 94 nsew signal output
rlabel metal2 s 95302 128302 95414 129102 6 io_out[25]
port 95 nsew signal output
rlabel metal3 s 0 14908 800 15148 6 io_out[26]
port 96 nsew signal output
rlabel metal2 s 99810 128302 99922 129102 6 io_out[27]
port 97 nsew signal output
rlabel metal2 s 44426 0 44538 800 6 io_out[28]
port 98 nsew signal output
rlabel metal3 s 127790 4028 128590 4268 6 io_out[29]
port 99 nsew signal output
rlabel metal2 s 18666 0 18778 800 6 io_out[2]
port 100 nsew signal output
rlabel metal3 s 0 16948 800 17188 6 io_out[30]
port 101 nsew signal output
rlabel metal3 s 0 37348 800 37588 6 io_out[31]
port 102 nsew signal output
rlabel metal3 s 0 122348 800 122588 6 io_out[32]
port 103 nsew signal output
rlabel metal3 s 127790 18988 128590 19228 6 io_out[33]
port 104 nsew signal output
rlabel metal3 s 127790 106028 128590 106268 6 io_out[34]
port 105 nsew signal output
rlabel metal3 s 127790 98548 128590 98788 6 io_out[35]
port 106 nsew signal output
rlabel metal2 s 40562 128302 40674 129102 6 io_out[36]
port 107 nsew signal output
rlabel metal3 s 127790 116228 128590 116468 6 io_out[37]
port 108 nsew signal output
rlabel metal3 s 0 112148 800 112388 6 io_out[3]
port 109 nsew signal output
rlabel metal3 s 127790 76108 128590 76348 6 io_out[4]
port 110 nsew signal output
rlabel metal2 s 59882 128302 59994 129102 6 io_out[5]
port 111 nsew signal output
rlabel metal2 s 123638 128302 123750 129102 6 io_out[6]
port 112 nsew signal output
rlabel metal3 s 0 52308 800 52548 6 io_out[7]
port 113 nsew signal output
rlabel metal2 s 49578 0 49690 800 6 io_out[8]
port 114 nsew signal output
rlabel metal3 s 0 39388 800 39628 6 io_out[9]
port 115 nsew signal output
rlabel metal3 s 127790 21028 128590 21268 6 la1_data_in[0]
port 116 nsew signal input
rlabel metal2 s 56662 0 56774 800 6 la1_data_in[10]
port 117 nsew signal input
rlabel metal3 s 127790 16268 128590 16508 6 la1_data_in[11]
port 118 nsew signal input
rlabel metal3 s 0 97188 800 97428 6 la1_data_in[12]
port 119 nsew signal input
rlabel metal2 s 87574 0 87686 800 6 la1_data_in[13]
port 120 nsew signal input
rlabel metal3 s 0 34628 800 34868 6 la1_data_in[14]
port 121 nsew signal input
rlabel metal2 s 43138 128302 43250 129102 6 la1_data_in[15]
port 122 nsew signal input
rlabel metal2 s 81134 128302 81246 129102 6 la1_data_in[16]
port 123 nsew signal input
rlabel metal2 s 61814 128302 61926 129102 6 la1_data_in[17]
port 124 nsew signal input
rlabel metal2 s 113334 0 113446 800 6 la1_data_in[18]
port 125 nsew signal input
rlabel metal2 s 45714 128302 45826 129102 6 la1_data_in[19]
port 126 nsew signal input
rlabel metal2 s 51510 0 51622 800 6 la1_data_in[1]
port 127 nsew signal input
rlabel metal3 s 0 94468 800 94708 6 la1_data_in[20]
port 128 nsew signal input
rlabel metal2 s 126214 128302 126326 129102 6 la1_data_in[21]
port 129 nsew signal input
rlabel metal3 s 127790 23748 128590 23988 6 la1_data_in[22]
port 130 nsew signal input
rlabel metal3 s 0 1988 800 2228 6 la1_data_in[23]
port 131 nsew signal input
rlabel metal2 s 37342 0 37454 800 6 la1_data_in[24]
port 132 nsew signal input
rlabel metal3 s 0 99908 800 100148 6 la1_data_in[25]
port 133 nsew signal input
rlabel metal3 s 127790 8788 128590 9028 6 la1_data_in[26]
port 134 nsew signal input
rlabel metal2 s 75338 0 75450 800 6 la1_data_in[27]
port 135 nsew signal input
rlabel metal3 s 0 86988 800 87228 6 la1_data_in[28]
port 136 nsew signal input
rlabel metal2 s 2566 128302 2678 129102 6 la1_data_in[29]
port 137 nsew signal input
rlabel metal2 s 30258 0 30370 800 6 la1_data_in[2]
port 138 nsew signal input
rlabel metal2 s 4498 0 4610 800 6 la1_data_in[30]
port 139 nsew signal input
rlabel metal2 s 99166 0 99278 800 6 la1_data_in[31]
port 140 nsew signal input
rlabel metal3 s 0 82228 800 82468 6 la1_data_in[3]
port 141 nsew signal input
rlabel metal2 s 109470 128302 109582 129102 6 la1_data_in[4]
port 142 nsew signal input
rlabel metal3 s 127790 63868 128590 64108 6 la1_data_in[5]
port 143 nsew signal input
rlabel metal2 s 50222 128302 50334 129102 6 la1_data_in[6]
port 144 nsew signal input
rlabel metal3 s 0 59788 800 60028 6 la1_data_in[7]
port 145 nsew signal input
rlabel metal2 s 52798 128302 52910 129102 6 la1_data_in[8]
port 146 nsew signal input
rlabel metal3 s 0 89708 800 89948 6 la1_data_in[9]
port 147 nsew signal input
rlabel metal2 s 21242 0 21354 800 6 la1_data_out[0]
port 148 nsew signal output
rlabel metal3 s 127790 31228 128590 31468 6 la1_data_out[10]
port 149 nsew signal output
rlabel metal2 s 58594 0 58706 800 6 la1_data_out[11]
port 150 nsew signal output
rlabel metal3 s 127790 118948 128590 119188 6 la1_data_out[12]
port 151 nsew signal output
rlabel metal2 s 12226 128302 12338 129102 6 la1_data_out[13]
port 152 nsew signal output
rlabel metal2 s 69542 128302 69654 129102 6 la1_data_out[14]
port 153 nsew signal output
rlabel metal3 s 0 4708 800 4948 6 la1_data_out[15]
port 154 nsew signal output
rlabel metal3 s 127790 43468 128590 43708 6 la1_data_out[16]
port 155 nsew signal output
rlabel metal3 s 127790 93788 128590 94028 6 la1_data_out[17]
port 156 nsew signal output
rlabel metal2 s 14802 128302 14914 129102 6 la1_data_out[18]
port 157 nsew signal output
rlabel metal3 s 127790 66588 128590 66828 6 la1_data_out[19]
port 158 nsew signal output
rlabel metal3 s 0 116908 800 117148 6 la1_data_out[1]
port 159 nsew signal output
rlabel metal3 s 0 27148 800 27388 6 la1_data_out[20]
port 160 nsew signal output
rlabel metal3 s 127790 111468 128590 111708 6 la1_data_out[21]
port 161 nsew signal output
rlabel metal2 s 78558 128302 78670 129102 6 la1_data_out[22]
port 162 nsew signal output
rlabel metal2 s 32834 0 32946 800 6 la1_data_out[23]
port 163 nsew signal output
rlabel metal3 s 127790 48908 128590 49148 6 la1_data_out[24]
port 164 nsew signal output
rlabel metal3 s 0 9468 800 9708 6 la1_data_out[25]
port 165 nsew signal output
rlabel metal3 s 127790 13548 128590 13788 6 la1_data_out[26]
port 166 nsew signal output
rlabel metal3 s 0 124388 800 124628 6 la1_data_out[27]
port 167 nsew signal output
rlabel metal2 s 115910 0 116022 800 6 la1_data_out[28]
port 168 nsew signal output
rlabel metal2 s 16090 0 16202 800 6 la1_data_out[29]
port 169 nsew signal output
rlabel metal2 s 54086 0 54198 800 6 la1_data_out[2]
port 170 nsew signal output
rlabel metal3 s 127790 33948 128590 34188 6 la1_data_out[30]
port 171 nsew signal output
rlabel metal3 s 127790 126428 128590 126668 6 la1_data_out[31]
port 172 nsew signal output
rlabel metal3 s 0 24428 800 24668 6 la1_data_out[3]
port 173 nsew signal output
rlabel metal2 s 117842 0 117954 800 6 la1_data_out[4]
port 174 nsew signal output
rlabel metal2 s 9006 0 9118 800 6 la1_data_out[5]
port 175 nsew signal output
rlabel metal3 s 127790 53668 128590 53908 6 la1_data_out[6]
port 176 nsew signal output
rlabel metal2 s 1922 0 2034 800 6 la1_data_out[7]
port 177 nsew signal output
rlabel metal3 s 127790 96508 128590 96748 6 la1_data_out[8]
port 178 nsew signal output
rlabel metal2 s 121062 128302 121174 129102 6 la1_data_out[9]
port 179 nsew signal output
rlabel metal2 s 127502 0 127614 800 6 la1_oenb[0]
port 180 nsew signal input
rlabel metal2 s 116554 128302 116666 129102 6 la1_oenb[10]
port 181 nsew signal input
rlabel metal3 s 0 72028 800 72268 6 la1_oenb[11]
port 182 nsew signal input
rlabel metal3 s 0 77468 800 77708 6 la1_oenb[12]
port 183 nsew signal input
rlabel metal2 s 77914 0 78026 800 6 la1_oenb[13]
port 184 nsew signal input
rlabel metal2 s -10 0 102 800 6 la1_oenb[14]
port 185 nsew signal input
rlabel metal2 s 92082 0 92194 800 6 la1_oenb[15]
port 186 nsew signal input
rlabel metal3 s 0 92428 800 92668 6 la1_oenb[16]
port 187 nsew signal input
rlabel metal2 s 10294 128302 10406 129102 6 la1_oenb[17]
port 188 nsew signal input
rlabel metal2 s 57306 128302 57418 129102 6 la1_oenb[18]
port 189 nsew signal input
rlabel metal3 s 0 69988 800 70228 6 la1_oenb[19]
port 190 nsew signal input
rlabel metal2 s 23174 0 23286 800 6 la1_oenb[1]
port 191 nsew signal input
rlabel metal2 s 7074 0 7186 800 6 la1_oenb[20]
port 192 nsew signal input
rlabel metal2 s 83710 128302 83822 129102 6 la1_oenb[21]
port 193 nsew signal input
rlabel metal2 s 54730 128302 54842 129102 6 la1_oenb[22]
port 194 nsew signal input
rlabel metal2 s 63746 0 63858 800 6 la1_oenb[23]
port 195 nsew signal input
rlabel metal2 s 102386 128302 102498 129102 6 la1_oenb[24]
port 196 nsew signal input
rlabel metal3 s 127790 26468 128590 26708 6 la1_oenb[25]
port 197 nsew signal input
rlabel metal3 s 0 101948 800 102188 6 la1_oenb[26]
port 198 nsew signal input
rlabel metal3 s 127790 91068 128590 91308 6 la1_oenb[27]
port 199 nsew signal input
rlabel metal2 s 25750 0 25862 800 6 la1_oenb[28]
port 200 nsew signal input
rlabel metal2 s 47002 0 47114 800 6 la1_oenb[29]
port 201 nsew signal input
rlabel metal3 s 0 22388 800 22628 6 la1_oenb[2]
port 202 nsew signal input
rlabel metal3 s 127790 89028 128590 89268 6 la1_oenb[30]
port 203 nsew signal input
rlabel metal2 s 73406 0 73518 800 6 la1_oenb[31]
port 204 nsew signal input
rlabel metal2 s 90794 128302 90906 129102 6 la1_oenb[3]
port 205 nsew signal input
rlabel metal2 s 88218 128302 88330 129102 6 la1_oenb[4]
port 206 nsew signal input
rlabel metal3 s 0 127108 800 127348 6 la1_oenb[5]
port 207 nsew signal input
rlabel metal2 s 19310 128302 19422 129102 6 la1_oenb[6]
port 208 nsew signal input
rlabel metal2 s 89506 0 89618 800 6 la1_oenb[7]
port 209 nsew signal input
rlabel metal3 s 0 31908 800 32148 6 la1_oenb[8]
port 210 nsew signal input
rlabel metal3 s 0 109428 800 109668 6 la1_oenb[9]
port 211 nsew signal input
rlabel metal4 s 4208 496 4528 126800 6 vccd1
port 212 nsew power input
rlabel metal4 s 34928 496 35248 126800 6 vccd1
port 212 nsew power input
rlabel metal4 s 65648 496 65968 126800 6 vccd1
port 212 nsew power input
rlabel metal4 s 96368 496 96688 126800 6 vccd1
port 212 nsew power input
rlabel metal4 s 19568 496 19888 126800 6 vssd1
port 213 nsew ground input
rlabel metal4 s 50288 496 50608 126800 6 vssd1
port 213 nsew ground input
rlabel metal4 s 81008 496 81328 126800 6 vssd1
port 213 nsew ground input
rlabel metal4 s 111728 496 112048 126800 6 vssd1
port 213 nsew ground input
rlabel metal3 s 127790 61148 128590 61388 6 wb_clk_i
port 214 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 128590 129102
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 35236652
string GDS_FILE /openlane/designs/wrapped_tetris/runs/RUN_2022.03.22_05.36.57/results/finishing/wrapped_tetris.magic.gds
string GDS_START 1432222
<< end >>

