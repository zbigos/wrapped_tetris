magic
tech sky130A
magscale 1 2
timestamp 1647922149
<< obsli1 >>
rect 1104 527 141312 140369
<< obsm1 >>
rect 14 496 142402 140400
<< metal2 >>
rect 3210 142181 3322 142981
rect 31546 142181 31658 142981
rect 59238 142181 59350 142981
rect 86930 142181 87042 142981
rect 114622 142181 114734 142981
rect 142314 142181 142426 142981
rect -10 0 102 800
rect 27682 0 27794 800
rect 55374 0 55486 800
rect 83066 0 83178 800
rect 110758 0 110870 800
rect 139094 0 139206 800
<< obsm2 >>
rect 20 142125 3154 142338
rect 3378 142125 31490 142338
rect 31714 142125 59182 142338
rect 59406 142125 86874 142338
rect 87098 142125 114566 142338
rect 114790 142125 142258 142338
rect 20 856 142396 142125
rect 158 496 27626 856
rect 27850 496 55318 856
rect 55542 496 83010 856
rect 83234 496 110702 856
rect 110926 496 139038 856
rect 139262 496 142396 856
<< metal3 >>
rect 0 116908 800 117148
rect 141669 112828 142469 113068
rect 0 87668 800 87908
rect 141669 83588 142469 83828
rect 0 58428 800 58668
rect 141669 54348 142469 54588
rect 0 29188 800 29428
rect 141669 25108 142469 25348
<< obsm3 >>
rect 800 117228 141669 140385
rect 880 116828 141669 117228
rect 800 113148 141669 116828
rect 800 112748 141589 113148
rect 800 87988 141669 112748
rect 880 87588 141669 87988
rect 800 83908 141669 87588
rect 800 83508 141589 83908
rect 800 58748 141669 83508
rect 880 58348 141669 58748
rect 800 54668 141669 58348
rect 800 54268 141589 54668
rect 800 29508 141669 54268
rect 880 29108 141669 29508
rect 800 25428 141669 29108
rect 800 25028 141589 25428
rect 800 511 141669 25028
<< metal4 >>
rect 4208 496 4528 140400
rect 19568 496 19888 140400
rect 34928 496 35248 140400
rect 50288 496 50608 140400
rect 65648 496 65968 140400
rect 81008 496 81328 140400
rect 96368 496 96688 140400
rect 111728 496 112048 140400
rect 127088 496 127408 140400
<< obsm4 >>
rect 4659 12411 19488 127125
rect 19968 12411 34848 127125
rect 35328 12411 50208 127125
rect 50688 12411 65568 127125
rect 66048 12411 80928 127125
rect 81408 12411 96288 127125
rect 96768 12411 103165 127125
<< labels >>
rlabel metal3 s 141669 25108 142469 25348 6 butt1
port 1 nsew signal input
rlabel metal2 s 142314 142181 142426 142981 6 butt2
port 2 nsew signal input
rlabel metal2 s 86930 142181 87042 142981 6 butt3
port 3 nsew signal input
rlabel metal2 s 55374 0 55486 800 6 butt4
port 4 nsew signal input
rlabel metal3 s 141669 112828 142469 113068 6 clk
port 5 nsew signal input
rlabel metal2 s 139094 0 139206 800 6 reset
port 6 nsew signal input
rlabel metal4 s 4208 496 4528 140400 6 vccd1
port 7 nsew power input
rlabel metal4 s 34928 496 35248 140400 6 vccd1
port 7 nsew power input
rlabel metal4 s 65648 496 65968 140400 6 vccd1
port 7 nsew power input
rlabel metal4 s 96368 496 96688 140400 6 vccd1
port 7 nsew power input
rlabel metal4 s 127088 496 127408 140400 6 vccd1
port 7 nsew power input
rlabel metal3 s 0 116908 800 117148 6 vga_b[0]
port 8 nsew signal output
rlabel metal2 s 59238 142181 59350 142981 6 vga_b[1]
port 9 nsew signal output
rlabel metal2 s -10 0 102 800 6 vga_b[2]
port 10 nsew signal output
rlabel metal2 s 31546 142181 31658 142981 6 vga_b[3]
port 11 nsew signal output
rlabel metal2 s 110758 0 110870 800 6 vga_g[0]
port 12 nsew signal output
rlabel metal2 s 27682 0 27794 800 6 vga_g[1]
port 13 nsew signal output
rlabel metal3 s 0 29188 800 29428 6 vga_g[2]
port 14 nsew signal output
rlabel metal3 s 141669 83588 142469 83828 6 vga_g[3]
port 15 nsew signal output
rlabel metal3 s 0 58428 800 58668 6 vga_h_sync
port 16 nsew signal output
rlabel metal2 s 114622 142181 114734 142981 6 vga_r[0]
port 17 nsew signal output
rlabel metal2 s 83066 0 83178 800 6 vga_r[1]
port 18 nsew signal output
rlabel metal3 s 0 87668 800 87908 6 vga_r[2]
port 19 nsew signal output
rlabel metal2 s 3210 142181 3322 142981 6 vga_r[3]
port 20 nsew signal output
rlabel metal3 s 141669 54348 142469 54588 6 vga_v_sync
port 21 nsew signal output
rlabel metal4 s 19568 496 19888 140400 6 vssd1
port 22 nsew ground input
rlabel metal4 s 50288 496 50608 140400 6 vssd1
port 22 nsew ground input
rlabel metal4 s 81008 496 81328 140400 6 vssd1
port 22 nsew ground input
rlabel metal4 s 111728 496 112048 140400 6 vssd1
port 22 nsew ground input
<< properties >>
string FIXED_BBOX 0 0 142469 142981
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 35409732
string GDS_FILE /openlane/designs/wrapped_tetris/runs/RUN_2022.03.22_04.02.55/results/finishing/top.magic.gds
string GDS_START 1399078
<< end >>

