* NGSPICE file created from wrapped_tetris.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_12 abstract view
.subckt sky130_fd_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_4 abstract view
.subckt sky130_fd_sc_hd__xor2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_2 abstract view
.subckt sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_1 abstract view
.subckt sky130_fd_sc_hd__mux4_1 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_4 abstract view
.subckt sky130_fd_sc_hd__or3b_4 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__ebufn_8 abstract view
.subckt sky130_fd_sc_hd__ebufn_8 A TE_B VGND VNB VPB VPWR Z
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_4 abstract view
.subckt sky130_fd_sc_hd__xnor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32oi_4 abstract view
.subckt sky130_fd_sc_hd__a32oi_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_2 abstract view
.subckt sky130_fd_sc_hd__a211oi_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_4 abstract view
.subckt sky130_fd_sc_hd__dfxtp_4 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_2 abstract view
.subckt sky130_fd_sc_hd__a221o_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_2 abstract view
.subckt sky130_fd_sc_hd__xor2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_2 abstract view
.subckt sky130_fd_sc_hd__nor3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_1 abstract view
.subckt sky130_fd_sc_hd__or2b_1 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_12 abstract view
.subckt sky130_fd_sc_hd__buf_12 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_2 abstract view
.subckt sky130_fd_sc_hd__mux4_2 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_1 abstract view
.subckt sky130_fd_sc_hd__o31ai_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_2 abstract view
.subckt sky130_fd_sc_hd__clkinv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_1 abstract view
.subckt sky130_fd_sc_hd__o22ai_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_1 abstract view
.subckt sky130_fd_sc_hd__o221ai_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_2 abstract view
.subckt sky130_fd_sc_hd__a41o_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_4 abstract view
.subckt sky130_fd_sc_hd__a21o_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_8 abstract view
.subckt sky130_fd_sc_hd__nor2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_2 abstract view
.subckt sky130_fd_sc_hd__and3b_2 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_1 abstract view
.subckt sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_1 abstract view
.subckt sky130_fd_sc_hd__nand4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_1 abstract view
.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_4 abstract view
.subckt sky130_fd_sc_hd__or4b_4 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_2 abstract view
.subckt sky130_fd_sc_hd__a211o_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_4 abstract view
.subckt sky130_fd_sc_hd__a221o_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_4 abstract view
.subckt sky130_fd_sc_hd__and2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_2 abstract view
.subckt sky130_fd_sc_hd__o21a_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_4 abstract view
.subckt sky130_fd_sc_hd__o211a_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_4 abstract view
.subckt sky130_fd_sc_hd__inv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_2 abstract view
.subckt sky130_fd_sc_hd__xnor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_2 abstract view
.subckt sky130_fd_sc_hd__nor4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_4 abstract view
.subckt sky130_fd_sc_hd__and3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_2 abstract view
.subckt sky130_fd_sc_hd__o31a_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311oi_1 abstract view
.subckt sky130_fd_sc_hd__a311oi_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_2 abstract view
.subckt sky130_fd_sc_hd__or4b_2 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_2 abstract view
.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_4 abstract view
.subckt sky130_fd_sc_hd__a21bo_4 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_2 abstract view
.subckt sky130_fd_sc_hd__nand2b_2 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_4 abstract view
.subckt sky130_fd_sc_hd__nand4_4 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_2 abstract view
.subckt sky130_fd_sc_hd__a31oi_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_2 abstract view
.subckt sky130_fd_sc_hd__nand3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111oi_1 abstract view
.subckt sky130_fd_sc_hd__a2111oi_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_2 abstract view
.subckt sky130_fd_sc_hd__a22oi_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_2 abstract view
.subckt sky130_fd_sc_hd__and2b_2 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_4 abstract view
.subckt sky130_fd_sc_hd__nor3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_4 abstract view
.subckt sky130_fd_sc_hd__nand2b_4 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_1 abstract view
.subckt sky130_fd_sc_hd__o41a_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_4 abstract view
.subckt sky130_fd_sc_hd__o221ai_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_2 abstract view
.subckt sky130_fd_sc_hd__a31o_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311ai_4 abstract view
.subckt sky130_fd_sc_hd__o311ai_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_4 abstract view
.subckt sky130_fd_sc_hd__o311a_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_4 abstract view
.subckt sky130_fd_sc_hd__nand3b_4 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4b_2 abstract view
.subckt sky130_fd_sc_hd__nor4b_2 A B C D_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_2 abstract view
.subckt sky130_fd_sc_hd__or2b_2 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_4 abstract view
.subckt sky130_fd_sc_hd__nor4_4 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_2 abstract view
.subckt sky130_fd_sc_hd__a21bo_2 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_1 abstract view
.subckt sky130_fd_sc_hd__a22oi_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_2 abstract view
.subckt sky130_fd_sc_hd__a311o_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_2 abstract view
.subckt sky130_fd_sc_hd__o2111ai_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_4 abstract view
.subckt sky130_fd_sc_hd__o31ai_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311ai_1 abstract view
.subckt sky130_fd_sc_hd__o311ai_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_2 abstract view
.subckt sky130_fd_sc_hd__o211a_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_2 abstract view
.subckt sky130_fd_sc_hd__o21bai_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_4 abstract view
.subckt sky130_fd_sc_hd__clkinv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_1 abstract view
.subckt sky130_fd_sc_hd__a31oi_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_4 abstract view
.subckt sky130_fd_sc_hd__and4bb_4 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_4 abstract view
.subckt sky130_fd_sc_hd__nand3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_2 abstract view
.subckt sky130_fd_sc_hd__o211ai_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_4 abstract view
.subckt sky130_fd_sc_hd__and4b_4 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_2 abstract view
.subckt sky130_fd_sc_hd__o32a_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_1 abstract view
.subckt sky130_fd_sc_hd__nand3b_1 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4b_4 abstract view
.subckt sky130_fd_sc_hd__nor4b_4 A B C D_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_2 abstract view
.subckt sky130_fd_sc_hd__a22o_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_4 abstract view
.subckt sky130_fd_sc_hd__and4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_4 abstract view
.subckt sky130_fd_sc_hd__and2b_4 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_4 abstract view
.subckt sky130_fd_sc_hd__o31a_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_1 abstract view
.subckt sky130_fd_sc_hd__a221oi_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_2 abstract view
.subckt sky130_fd_sc_hd__a21o_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_1 abstract view
.subckt sky130_fd_sc_hd__nor3b_1 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41oi_1 abstract view
.subckt sky130_fd_sc_hd__a41oi_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_2 abstract view
.subckt sky130_fd_sc_hd__nand3b_2 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_4 abstract view
.subckt sky130_fd_sc_hd__a22oi_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkdlybuf4s25_1 abstract view
.subckt sky130_fd_sc_hd__clkdlybuf4s25_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_2 abstract view
.subckt sky130_fd_sc_hd__or3b_2 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_4 abstract view
.subckt sky130_fd_sc_hd__a21boi_4 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkdlybuf4s50_1 abstract view
.subckt sky130_fd_sc_hd__clkdlybuf4s50_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_2 abstract view
.subckt sky130_fd_sc_hd__nor3b_2 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_2 abstract view
.subckt sky130_fd_sc_hd__o21ba_2 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_4 abstract view
.subckt sky130_fd_sc_hd__nor3b_4 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_4 abstract view
.subckt sky130_fd_sc_hd__a2111o_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2b_2 abstract view
.subckt sky130_fd_sc_hd__nor2b_2 A B_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2b_4 abstract view
.subckt sky130_fd_sc_hd__nor2b_4 A B_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_8 abstract view
.subckt sky130_fd_sc_hd__nand2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_2 abstract view
.subckt sky130_fd_sc_hd__a32o_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_4 abstract view
.subckt sky130_fd_sc_hd__or4bb_4 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_2 abstract view
.subckt sky130_fd_sc_hd__or4bb_2 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_2 abstract view
.subckt sky130_fd_sc_hd__o311a_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_2 abstract view
.subckt sky130_fd_sc_hd__o22ai_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_4 abstract view
.subckt sky130_fd_sc_hd__o211ai_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_2 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_4 abstract view
.subckt sky130_fd_sc_hd__a31oi_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311oi_2 abstract view
.subckt sky130_fd_sc_hd__a311oi_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_2 abstract view
.subckt sky130_fd_sc_hd__a2111o_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_4 abstract view
.subckt sky130_fd_sc_hd__mux2_4 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_4 abstract view
.subckt sky130_fd_sc_hd__and3b_4 A_N B C VGND VNB VPB VPWR X
.ends

.subckt wrapped_tetris active io_in[0] io_in[10] io_in[11] io_in[12] io_in[13] io_in[14]
+ io_in[15] io_in[16] io_in[17] io_in[18] io_in[19] io_in[1] io_in[20] io_in[21] io_in[22]
+ io_in[23] io_in[24] io_in[25] io_in[26] io_in[27] io_in[28] io_in[29] io_in[2] io_in[30]
+ io_in[31] io_in[32] io_in[33] io_in[34] io_in[35] io_in[36] io_in[37] io_in[3] io_in[4]
+ io_in[5] io_in[6] io_in[7] io_in[8] io_in[9] io_oeb[0] io_oeb[10] io_oeb[11] io_oeb[12]
+ io_oeb[13] io_oeb[14] io_oeb[15] io_oeb[16] io_oeb[17] io_oeb[18] io_oeb[19] io_oeb[1]
+ io_oeb[20] io_oeb[21] io_oeb[22] io_oeb[23] io_oeb[24] io_oeb[25] io_oeb[26] io_oeb[27]
+ io_oeb[28] io_oeb[29] io_oeb[2] io_oeb[30] io_oeb[31] io_oeb[32] io_oeb[33] io_oeb[34]
+ io_oeb[35] io_oeb[36] io_oeb[37] io_oeb[3] io_oeb[4] io_oeb[5] io_oeb[6] io_oeb[7]
+ io_oeb[8] io_oeb[9] io_out[0] io_out[10] io_out[11] io_out[12] io_out[13] io_out[14]
+ io_out[15] io_out[16] io_out[17] io_out[18] io_out[19] io_out[1] io_out[20] io_out[21]
+ io_out[22] io_out[23] io_out[24] io_out[25] io_out[26] io_out[27] io_out[28] io_out[29]
+ io_out[2] io_out[30] io_out[31] io_out[32] io_out[33] io_out[34] io_out[35] io_out[36]
+ io_out[37] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7] io_out[8] io_out[9]
+ la1_data_in[0] la1_data_in[10] la1_data_in[11] la1_data_in[12] la1_data_in[13] la1_data_in[14]
+ la1_data_in[15] la1_data_in[16] la1_data_in[17] la1_data_in[18] la1_data_in[19]
+ la1_data_in[1] la1_data_in[20] la1_data_in[21] la1_data_in[22] la1_data_in[23] la1_data_in[24]
+ la1_data_in[25] la1_data_in[26] la1_data_in[27] la1_data_in[28] la1_data_in[29]
+ la1_data_in[2] la1_data_in[30] la1_data_in[31] la1_data_in[3] la1_data_in[4] la1_data_in[5]
+ la1_data_in[6] la1_data_in[7] la1_data_in[8] la1_data_in[9] la1_data_out[0] la1_data_out[10]
+ la1_data_out[11] la1_data_out[12] la1_data_out[13] la1_data_out[14] la1_data_out[15]
+ la1_data_out[16] la1_data_out[17] la1_data_out[18] la1_data_out[19] la1_data_out[1]
+ la1_data_out[20] la1_data_out[21] la1_data_out[22] la1_data_out[23] la1_data_out[24]
+ la1_data_out[25] la1_data_out[26] la1_data_out[27] la1_data_out[28] la1_data_out[29]
+ la1_data_out[2] la1_data_out[30] la1_data_out[31] la1_data_out[3] la1_data_out[4]
+ la1_data_out[5] la1_data_out[6] la1_data_out[7] la1_data_out[8] la1_data_out[9]
+ la1_oenb[0] la1_oenb[10] la1_oenb[11] la1_oenb[12] la1_oenb[13] la1_oenb[14] la1_oenb[15]
+ la1_oenb[16] la1_oenb[17] la1_oenb[18] la1_oenb[19] la1_oenb[1] la1_oenb[20] la1_oenb[21]
+ la1_oenb[22] la1_oenb[23] la1_oenb[24] la1_oenb[25] la1_oenb[26] la1_oenb[27] la1_oenb[28]
+ la1_oenb[29] la1_oenb[2] la1_oenb[30] la1_oenb[31] la1_oenb[3] la1_oenb[4] la1_oenb[5]
+ la1_oenb[6] la1_oenb[7] la1_oenb[8] la1_oenb[9] vccd1 vssd1 wb_clk_i
XFILLER_228_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_227_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_223_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09671_ _12070_/A _12070_/B vssd1 vssd1 vccd1 vccd1 _09719_/B sky130_fd_sc_hd__xor2_4
XFILLER_80_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_1298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18869_ _18870_/CLK _18869_/D vssd1 vssd1 vccd1 vccd1 _18869_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_227_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_223_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XINSDIODE2_260 _13848_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_271 _18397_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_206_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09105_ _18740_/Q _18739_/Q _18738_/Q vssd1 vssd1 vccd1 vccd1 _09109_/A sky130_fd_sc_hd__or3_4
XFILLER_148_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_175_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09036_ _09040_/A vssd1 vssd1 vccd1 vccd1 _09036_/Y sky130_fd_sc_hd__inv_2
XFILLER_108_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_136_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_213_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09938_ _09413_/A _09408_/C _09418_/D _10956_/A _09937_/X _09909_/X vssd1 vssd1 vccd1
+ vccd1 _09938_/X sky130_fd_sc_hd__mux4_1
XFILLER_104_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_213_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09869_ _18107_/Q vssd1 vssd1 vccd1 vccd1 _09872_/A sky130_fd_sc_hd__inv_2
XFILLER_73_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11900_ _17793_/Q vssd1 vssd1 vccd1 vccd1 _12021_/A sky130_fd_sc_hd__inv_2
XTAP_3224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12880_ _12880_/A vssd1 vssd1 vccd1 vccd1 _17956_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_172_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11831_ _11591_/B _11830_/X _11899_/C vssd1 vssd1 vccd1 vccd1 _11832_/C sky130_fd_sc_hd__a21oi_1
XTAP_2534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14550_ _17602_/A _17635_/A vssd1 vssd1 vccd1 vccd1 _16817_/A sky130_fd_sc_hd__or2_4
XTAP_2578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11762_ _11767_/C _12509_/A _11767_/B vssd1 vssd1 vccd1 vccd1 _11763_/C sky130_fd_sc_hd__a21o_1
XTAP_1844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13501_ _13501_/A _17804_/Q _13518_/A vssd1 vssd1 vccd1 vccd1 _13557_/B sky130_fd_sc_hd__or3b_4
XFILLER_183_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10713_ _10770_/A vssd1 vssd1 vccd1 vccd1 _10743_/A sky130_fd_sc_hd__clkbuf_2
XTAP_1877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14481_ _14481_/A vssd1 vssd1 vccd1 vccd1 _18215_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11693_ _17850_/Q vssd1 vssd1 vccd1 vccd1 _11704_/C sky130_fd_sc_hd__clkbuf_2
XTAP_1899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16220_ _17410_/A _16366_/B vssd1 vssd1 vccd1 vccd1 _16289_/A sky130_fd_sc_hd__or2_1
XFILLER_224_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13432_ _13635_/A _13693_/A _13710_/C vssd1 vssd1 vccd1 vccd1 _13438_/B sky130_fd_sc_hd__a21oi_1
X_10644_ _10644_/A vssd1 vssd1 vccd1 vccd1 _10680_/A sky130_fd_sc_hd__buf_6
XFILLER_201_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16151_ _16173_/A vssd1 vssd1 vccd1 vccd1 _16170_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_167_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_220_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10575_ _10575_/A _10575_/B vssd1 vssd1 vccd1 vccd1 _10575_/X sky130_fd_sc_hd__or2_1
X_13363_ _14384_/B _13363_/B vssd1 vssd1 vccd1 vccd1 _13363_/Y sky130_fd_sc_hd__nand2_1
X_15102_ _15207_/A vssd1 vssd1 vccd1 vccd1 _15187_/A sky130_fd_sc_hd__clkbuf_2
X_12314_ _12314_/A vssd1 vssd1 vccd1 vccd1 _17879_/D sky130_fd_sc_hd__clkbuf_1
X_16082_ _16132_/A _16082_/B vssd1 vssd1 vccd1 vccd1 _16082_/Y sky130_fd_sc_hd__nand2_1
X_13294_ _18058_/Q _18061_/Q _18060_/Q _18063_/Q vssd1 vssd1 vccd1 vccd1 _13297_/A
+ sky130_fd_sc_hd__or4_1
XFILLER_177_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_182_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_170_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15033_ _18382_/Q _18346_/Q _15033_/S vssd1 vssd1 vccd1 vccd1 _15033_/X sky130_fd_sc_hd__mux2_1
XFILLER_68_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12245_ _17863_/Q _17860_/Q _12242_/X vssd1 vssd1 vccd1 vccd1 _12269_/C sky130_fd_sc_hd__a21o_1
XFILLER_181_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_1333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12176_ _12174_/X _12175_/Y _12163_/X vssd1 vssd1 vccd1 vccd1 _17846_/D sky130_fd_sc_hd__o21a_1
XFILLER_174_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11127_ _11455_/C vssd1 vssd1 vccd1 vccd1 _13446_/A sky130_fd_sc_hd__buf_2
XFILLER_228_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16984_ _16975_/A _17028_/C _18809_/Q vssd1 vssd1 vccd1 vccd1 _16984_/Y sky130_fd_sc_hd__o21bai_1
XFILLER_7_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15935_ _15984_/A _15935_/B _15964_/C vssd1 vssd1 vccd1 vccd1 _15935_/X sky130_fd_sc_hd__or3_1
X_18723_ _18724_/CLK _18723_/D vssd1 vssd1 vccd1 vccd1 _18723_/Q sky130_fd_sc_hd__dfxtp_2
X_11058_ _13448_/A _17816_/Q _12272_/A vssd1 vssd1 vccd1 vccd1 _11059_/A sky130_fd_sc_hd__mux2_1
XFILLER_49_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_60_wb_clk_i _18759_/CLK vssd1 vssd1 vccd1 vccd1 _18724_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_64_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10009_ _10009_/A vssd1 vssd1 vccd1 vccd1 _10010_/A sky130_fd_sc_hd__clkbuf_2
X_18654_ _18663_/CLK _18654_/D vssd1 vssd1 vccd1 vccd1 _18654_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_36_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15866_ _15865_/B _15864_/X _15865_/Y _15861_/X vssd1 vssd1 vccd1 vccd1 _18545_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_4470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14817_ _18330_/Q _18294_/Q _14830_/S vssd1 vssd1 vccd1 vccd1 _14817_/X sky130_fd_sc_hd__mux2_1
X_17605_ _17602_/Y _17604_/X _17591_/X vssd1 vssd1 vccd1 vccd1 _17605_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_91_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18585_ _18590_/CLK _18585_/D vssd1 vssd1 vccd1 vccd1 _18585_/Q sky130_fd_sc_hd__dfxtp_1
X_15797_ _15944_/A _15844_/B vssd1 vssd1 vccd1 vccd1 _15806_/B sky130_fd_sc_hd__nor2_1
XTAP_3780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17536_ _17536_/A _17536_/B vssd1 vssd1 vccd1 vccd1 _17544_/B sky130_fd_sc_hd__nor2_2
X_14748_ _14753_/B _14745_/X _14747_/X _14738_/X vssd1 vssd1 vccd1 vccd1 _18276_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_33_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_178_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_225_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17467_ _18965_/Q _18929_/Q _17467_/S vssd1 vssd1 vccd1 vccd1 _17467_/X sky130_fd_sc_hd__mux2_1
X_14679_ _14734_/A _14690_/B _15268_/B vssd1 vssd1 vccd1 vccd1 _14679_/X sky130_fd_sc_hd__or3_1
XFILLER_60_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_1359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_203_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16418_ _16456_/A vssd1 vssd1 vccd1 vccd1 _16418_/X sky130_fd_sc_hd__clkbuf_2
X_19206_ _19206_/A _08975_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[6] sky130_fd_sc_hd__ebufn_8
XFILLER_220_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17398_ _18948_/Q _18912_/Q _17406_/S vssd1 vssd1 vccd1 vccd1 _17398_/X sky130_fd_sc_hd__mux2_1
XFILLER_160_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_186_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_201_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19137_ _19137_/A _09042_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[7] sky130_fd_sc_hd__ebufn_8
X_16349_ _18694_/Q _18658_/Q _16363_/S vssd1 vssd1 vccd1 vccd1 _16349_/X sky130_fd_sc_hd__mux2_1
XFILLER_160_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_1367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_146_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_195_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_218_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18019_ _18095_/CLK _18019_/D vssd1 vssd1 vccd1 vccd1 _18019_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_161_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09723_ _09723_/A _09723_/B vssd1 vssd1 vccd1 vccd1 _10070_/B sky130_fd_sc_hd__xnor2_4
XFILLER_74_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09654_ _09692_/A _09654_/B vssd1 vssd1 vccd1 vccd1 _10582_/S sky130_fd_sc_hd__or2_4
XFILLER_82_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_216_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_215_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09585_ _09585_/A _09585_/B _09585_/C vssd1 vssd1 vccd1 vccd1 _09586_/B sky130_fd_sc_hd__or3_1
XTAP_1107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_230_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_204_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_1300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10360_ _10342_/X _10358_/X _10605_/C vssd1 vssd1 vccd1 vccd1 _10360_/X sky130_fd_sc_hd__o21a_1
XFILLER_124_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09019_ _09022_/A vssd1 vssd1 vccd1 vccd1 _09019_/Y sky130_fd_sc_hd__inv_2
XFILLER_151_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10291_ _10291_/A vssd1 vssd1 vccd1 vccd1 _10291_/X sky130_fd_sc_hd__buf_4
X_12030_ _12099_/B vssd1 vssd1 vccd1 vccd1 _13420_/A sky130_fd_sc_hd__buf_2
XFILLER_120_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13981_ _18343_/Q _13677_/X _13623_/A _18349_/Q vssd1 vssd1 vccd1 vccd1 _13981_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_63_1293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_219_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15720_ _15720_/A vssd1 vssd1 vccd1 vccd1 _15720_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_101_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12932_ _17993_/Q _12955_/A _12962_/A _11044_/B vssd1 vssd1 vccd1 vccd1 _12933_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_218_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19041__12 vssd1 vssd1 vccd1 vccd1 _19041__12/HI _19135_/A sky130_fd_sc_hd__conb_1
XTAP_3054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15651_ _15694_/A _15651_/B vssd1 vssd1 vccd1 vccd1 _15651_/Y sky130_fd_sc_hd__nand2_1
XFILLER_218_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12863_ _17951_/Q _12865_/C _12862_/X vssd1 vssd1 vccd1 vccd1 _12864_/B sky130_fd_sc_hd__o21ai_1
XTAP_3065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14602_ _14665_/A _14665_/B _15199_/B vssd1 vssd1 vccd1 vccd1 _14602_/X sky130_fd_sc_hd__or3_1
XTAP_2353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18370_ _18373_/CLK _18370_/D vssd1 vssd1 vccd1 vccd1 _18370_/Q sky130_fd_sc_hd__dfxtp_2
X_11814_ _17661_/A vssd1 vssd1 vccd1 vccd1 _17420_/A sky130_fd_sc_hd__buf_4
XTAP_2364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15582_ _15582_/A vssd1 vssd1 vccd1 vccd1 _15633_/A sky130_fd_sc_hd__clkbuf_2
XTAP_1630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12794_ _12646_/A _12792_/X _12646_/B _12793_/Y vssd1 vssd1 vccd1 vccd1 _12794_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_109_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_221_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_202_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_199_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17321_ _18928_/Q _18892_/Q _17347_/S vssd1 vssd1 vccd1 vccd1 _17321_/X sky130_fd_sc_hd__mux2_1
XFILLER_14_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14533_ _14533_/A vssd1 vssd1 vccd1 vccd1 _14533_/X sky130_fd_sc_hd__clkbuf_4
X_11745_ _11824_/A _11826_/C _11826_/B vssd1 vssd1 vccd1 vccd1 _11856_/A sky130_fd_sc_hd__a21o_1
XFILLER_42_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_5_29_0_wb_clk_i clkbuf_5_29_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_5_29_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_159_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17252_ _17275_/A _17252_/B vssd1 vssd1 vccd1 vccd1 _17252_/Y sky130_fd_sc_hd__nand2_1
XFILLER_53_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14464_ _14464_/A _14464_/B vssd1 vssd1 vccd1 vccd1 _14470_/C sky130_fd_sc_hd__and2_1
X_11676_ _11651_/A _11675_/Y _11848_/B _11640_/Y vssd1 vssd1 vccd1 vccd1 _11676_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_30_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16203_ _16202_/B _16201_/X _16202_/Y _16185_/X vssd1 vssd1 vccd1 vccd1 _18623_/D
+ sky130_fd_sc_hd__o211a_1
X_13415_ _13415_/A _13415_/B vssd1 vssd1 vccd1 vccd1 _13415_/Y sky130_fd_sc_hd__nor2_1
XFILLER_179_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17183_ _17471_/A _17256_/C vssd1 vssd1 vccd1 vccd1 _17189_/B sky130_fd_sc_hd__nor2_2
X_10627_ _18130_/Q _10627_/B vssd1 vssd1 vccd1 vccd1 _10656_/B sky130_fd_sc_hd__xnor2_4
X_14395_ _17564_/A _14395_/B vssd1 vssd1 vccd1 vccd1 _14396_/A sky130_fd_sc_hd__and2_1
XFILLER_183_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16134_ _16886_/A vssd1 vssd1 vccd1 vccd1 _16734_/A sky130_fd_sc_hd__buf_6
XFILLER_128_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13346_ _13346_/A vssd1 vssd1 vccd1 vccd1 _13346_/X sky130_fd_sc_hd__buf_2
XFILLER_154_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10558_ _10183_/A _10549_/X _10553_/X _10555_/X _10557_/X vssd1 vssd1 vccd1 vccd1
+ _10558_/Y sky130_fd_sc_hd__a32oi_4
XFILLER_182_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16065_ _18593_/Q _16064_/B _16064_/Y _16048_/X vssd1 vssd1 vccd1 vccd1 _18593_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_185_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13277_ _19010_/Q _19009_/Q _19012_/Q _19011_/Q vssd1 vssd1 vccd1 vccd1 _13278_/D
+ sky130_fd_sc_hd__or4_1
XFILLER_6_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10489_ _09148_/C _10722_/A _10489_/S vssd1 vssd1 vccd1 vccd1 _10489_/X sky130_fd_sc_hd__mux2_1
X_15016_ _15125_/A vssd1 vssd1 vccd1 vccd1 _15105_/A sky130_fd_sc_hd__buf_2
X_12228_ _11603_/A _12221_/A _12233_/C _12222_/X vssd1 vssd1 vccd1 vccd1 _12228_/Y
+ sky130_fd_sc_hd__a211oi_2
XFILLER_9_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12159_ _13458_/A vssd1 vssd1 vccd1 vccd1 _12172_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_151_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16967_ _17164_/A vssd1 vssd1 vccd1 vccd1 _17032_/A sky130_fd_sc_hd__buf_2
XFILLER_110_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18706_ _18708_/CLK _18706_/D vssd1 vssd1 vccd1 vccd1 _18706_/Q sky130_fd_sc_hd__dfxtp_2
X_15918_ _16034_/A vssd1 vssd1 vccd1 vccd1 _16014_/A sky130_fd_sc_hd__buf_2
X_16898_ _16954_/A _16903_/B vssd1 vssd1 vccd1 vccd1 _16898_/Y sky130_fd_sc_hd__nand2_1
XFILLER_65_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18637_ _18641_/CLK _18637_/D vssd1 vssd1 vccd1 vccd1 _18637_/Q sky130_fd_sc_hd__dfxtp_2
X_15849_ _18577_/Q _18541_/Q _15859_/S vssd1 vssd1 vccd1 vccd1 _15849_/X sky130_fd_sc_hd__mux2_1
XFILLER_25_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_212_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09370_ _09370_/A _09370_/B _09370_/C _10883_/A vssd1 vssd1 vccd1 vccd1 _09371_/C
+ sky130_fd_sc_hd__and4_1
X_18568_ _18607_/CLK _18568_/D vssd1 vssd1 vccd1 vccd1 _18568_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_75_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_224_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_206_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_221_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_220_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_177_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17519_ _17519_/A vssd1 vssd1 vccd1 vccd1 _17533_/S sky130_fd_sc_hd__clkbuf_2
X_18499_ _18504_/CLK _18499_/D vssd1 vssd1 vccd1 vccd1 _18499_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_127_1243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_177_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_178_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_229_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_134_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_4 _09058_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09706_ _10060_/A vssd1 vssd1 vccd1 vccd1 _10102_/S sky130_fd_sc_hd__buf_4
XFILLER_74_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09637_ _09637_/A _09637_/B vssd1 vssd1 vccd1 vccd1 _09637_/X sky130_fd_sc_hd__or2_1
XFILLER_3_1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_204_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_128_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_215_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09568_ _09568_/A vssd1 vssd1 vccd1 vccd1 _09600_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_93_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_212_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09499_ _18197_/Q _09499_/B vssd1 vssd1 vccd1 vccd1 _09500_/B sky130_fd_sc_hd__or2_1
XFILLER_230_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11530_ _11530_/A _11530_/B vssd1 vssd1 vccd1 vccd1 _11530_/X sky130_fd_sc_hd__and2_1
XFILLER_184_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_221_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11461_ _17885_/Q vssd1 vssd1 vccd1 vccd1 _11463_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_109_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13200_ _13208_/A _18057_/Q vssd1 vssd1 vccd1 vccd1 _13201_/A sky130_fd_sc_hd__and2_1
XFILLER_104_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10412_ _10412_/A vssd1 vssd1 vccd1 vccd1 _10413_/A sky130_fd_sc_hd__clkbuf_8
X_14180_ _18674_/Q _13515_/X _13546_/X _18671_/Q _14179_/X vssd1 vssd1 vccd1 vccd1
+ _14180_/X sky130_fd_sc_hd__a221o_1
XFILLER_136_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11392_ _13485_/A _11392_/B vssd1 vssd1 vccd1 vccd1 _11539_/B sky130_fd_sc_hd__nor2_1
XFILLER_165_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13131_ _13142_/A vssd1 vssd1 vccd1 vccd1 _13140_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_151_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10343_ _09126_/A _09136_/B _09131_/A _09126_/D _10274_/S _09905_/X vssd1 vssd1 vccd1
+ vccd1 _10343_/X sky130_fd_sc_hd__mux4_1
XFILLER_174_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_180_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10274_ _09160_/A _09165_/C _10274_/S vssd1 vssd1 vccd1 vccd1 _10274_/X sky130_fd_sc_hd__mux2_1
X_13062_ _18005_/Q _13082_/A _13085_/A vssd1 vssd1 vccd1 vccd1 _13063_/B sky130_fd_sc_hd__a21boi_1
XFILLER_65_1333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12013_ _12023_/B _11971_/B _13426_/A _11963_/A vssd1 vssd1 vccd1 vccd1 _12016_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_65_1366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17870_ _19030_/CLK _17870_/D vssd1 vssd1 vccd1 vccd1 _17870_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_61_1208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16821_ _16928_/A vssd1 vssd1 vccd1 vccd1 _16842_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_171_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16752_ _16752_/A _16755_/B vssd1 vssd1 vccd1 vccd1 _16752_/Y sky130_fd_sc_hd__nand2_1
XFILLER_4_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13964_ _18427_/Q _13580_/A _13734_/X _18421_/Q _13963_/X vssd1 vssd1 vccd1 vccd1
+ _13964_/X sky130_fd_sc_hd__a221o_1
XFILLER_219_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15703_ _15885_/A vssd1 vssd1 vccd1 vccd1 _15751_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_185_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12915_ _12913_/X _12915_/B _12915_/C vssd1 vssd1 vccd1 vccd1 _12916_/A sky130_fd_sc_hd__and3b_1
X_16683_ _16760_/A vssd1 vssd1 vccd1 vccd1 _16683_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13895_ _18622_/Q _13657_/A _13893_/X _13894_/X vssd1 vssd1 vccd1 vccd1 _13895_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_34_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18422_ _18423_/CLK _18422_/D vssd1 vssd1 vccd1 vccd1 _18422_/Q sky130_fd_sc_hd__dfxtp_4
X_15634_ _15633_/B _15632_/X _15633_/Y _15616_/X vssd1 vssd1 vccd1 vccd1 _18488_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_2150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12846_ _12846_/A _12846_/B vssd1 vssd1 vccd1 vccd1 _12848_/B sky130_fd_sc_hd__nand2_1
XFILLER_181_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18353_ _18356_/CLK _18353_/D vssd1 vssd1 vccd1 vccd1 _18353_/Q sky130_fd_sc_hd__dfxtp_4
XTAP_2194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15565_ _18508_/Q _18472_/Q _15565_/S vssd1 vssd1 vccd1 vccd1 _15565_/X sky130_fd_sc_hd__mux2_1
XFILLER_159_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12777_ _18002_/Q vssd1 vssd1 vccd1 vccd1 _13080_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_14_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17304_ _17304_/A vssd1 vssd1 vccd1 vccd1 _17304_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_1493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14516_ _14515_/B _14513_/B _18229_/Q vssd1 vssd1 vccd1 vccd1 _14516_/X sky130_fd_sc_hd__o21a_1
XFILLER_175_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18284_ _18290_/CLK _18284_/D vssd1 vssd1 vccd1 vccd1 _18284_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_9_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11728_ _11727_/Y _11727_/A _17915_/Q vssd1 vssd1 vccd1 vccd1 _11729_/S sky130_fd_sc_hd__mux2_1
XFILLER_230_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_226_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15496_ _15516_/A vssd1 vssd1 vccd1 vccd1 _15496_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_175_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17235_ _17240_/B _17233_/X _17234_/X _17219_/X vssd1 vssd1 vccd1 vccd1 _18870_/D
+ sky130_fd_sc_hd__o211a_1
X_14447_ _14445_/Y _14386_/Y _14446_/X _18202_/Q vssd1 vssd1 vccd1 vccd1 _14448_/B
+ sky130_fd_sc_hd__a22o_1
X_11659_ _11497_/B _11669_/A _11681_/C _11659_/D vssd1 vssd1 vccd1 vccd1 _11705_/D
+ sky130_fd_sc_hd__and4b_1
XFILLER_70_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17166_ _17169_/B _17163_/X _17165_/Y _17161_/X vssd1 vssd1 vccd1 vccd1 _18853_/D
+ sky130_fd_sc_hd__o211a_1
X_14378_ _14375_/X _14376_/Y _17766_/A vssd1 vssd1 vccd1 vccd1 _18187_/D sky130_fd_sc_hd__a21oi_1
XFILLER_128_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16117_ _16173_/A vssd1 vssd1 vccd1 vccd1 _16145_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_116_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13329_ _18093_/Q _13329_/B _13314_/A vssd1 vssd1 vccd1 vccd1 _13329_/X sky130_fd_sc_hd__or3b_1
XFILLER_192_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17097_ _17105_/B _17094_/X _17095_/X _17096_/X vssd1 vssd1 vccd1 vccd1 _18837_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_50_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16048_ _16139_/A vssd1 vssd1 vccd1 vccd1 _16048_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_192_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_215_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_229_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17999_ _18997_/CLK _17999_/D vssd1 vssd1 vccd1 vccd1 _17999_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_56_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_226_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_1310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_226_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09422_ _09427_/B _09450_/A _09420_/X _09421_/Y vssd1 vssd1 vccd1 vccd1 _09423_/B
+ sky130_fd_sc_hd__o31a_1
XFILLER_44_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09353_ _18443_/Q _18442_/Q _18441_/Q vssd1 vssd1 vccd1 vccd1 _09354_/D sky130_fd_sc_hd__or3_4
XFILLER_40_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09284_ _18872_/Q _18871_/Q _18870_/Q vssd1 vssd1 vccd1 vccd1 _09287_/B sky130_fd_sc_hd__or3_4
XFILLER_166_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_1232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_193_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_175_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_173_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_216_1366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08999_ _09003_/A vssd1 vssd1 vccd1 vccd1 _08999_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_188_wb_clk_i clkbuf_5_9_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17890_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_134_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_229_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_1274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_216_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_117_wb_clk_i clkbuf_5_30_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18485_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_28_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10961_ _09365_/A _09370_/B _10883_/A _09360_/C _10003_/S _10017_/S vssd1 vssd1 vccd1
+ vccd1 _10962_/B sky130_fd_sc_hd__mux4_1
XFILLER_95_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12700_ _12699_/Y _12691_/B _17934_/Q vssd1 vssd1 vccd1 vccd1 _12700_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_216_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13680_ _18543_/Q _13529_/A _13535_/A _18519_/Q vssd1 vssd1 vccd1 vccd1 _13680_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_3_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10892_ _09386_/A _09376_/B _09381_/C _09972_/A _10060_/A _10025_/A vssd1 vssd1 vccd1
+ vccd1 _10892_/X sky130_fd_sc_hd__mux4_1
XFILLER_182_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12631_ _12618_/A _12619_/A _12618_/B _12630_/X vssd1 vssd1 vccd1 vccd1 _12632_/B
+ sky130_fd_sc_hd__o31a_1
XFILLER_34_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15350_ _15352_/B _15348_/X _15349_/Y _15340_/X vssd1 vssd1 vccd1 vccd1 _18421_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_70_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_223_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12562_ _17923_/Q vssd1 vssd1 vccd1 vccd1 _12594_/B sky130_fd_sc_hd__inv_2
XFILLER_184_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_212_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_197_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14301_ _18176_/Q vssd1 vssd1 vccd1 vccd1 _15463_/B sky130_fd_sc_hd__buf_2
XFILLER_106_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_211_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11513_ _11513_/A _11534_/A vssd1 vssd1 vccd1 vccd1 _11513_/Y sky130_fd_sc_hd__nand2_1
X_15281_ _18445_/Q _18409_/Q _15285_/S vssd1 vssd1 vccd1 vccd1 _15281_/X sky130_fd_sc_hd__mux2_1
XFILLER_11_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12493_ _17910_/Q _12493_/B vssd1 vssd1 vccd1 vccd1 _12495_/D sky130_fd_sc_hd__xor2_1
XFILLER_221_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17020_ _17096_/A vssd1 vssd1 vccd1 vccd1 _17020_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_8_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14232_ _14202_/X _14226_/Y _14231_/X _13334_/X vssd1 vssd1 vccd1 vccd1 _18169_/D
+ sky130_fd_sc_hd__o211a_1
X_11444_ _11438_/X _11441_/Y _11443_/X vssd1 vssd1 vccd1 vccd1 _11444_/X sky130_fd_sc_hd__o21a_1
XFILLER_32_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14163_ _18971_/Q _14124_/X _13538_/A _18953_/Q vssd1 vssd1 vccd1 vccd1 _14163_/X
+ sky130_fd_sc_hd__a22o_1
X_11375_ _11375_/A _11375_/B vssd1 vssd1 vccd1 vccd1 _11376_/B sky130_fd_sc_hd__or2_1
XFILLER_124_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13114_ _13118_/A _18018_/Q vssd1 vssd1 vccd1 vccd1 _13115_/A sky130_fd_sc_hd__and2_1
XFILLER_180_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10326_ _10324_/X _10325_/X _10333_/S vssd1 vssd1 vccd1 vccd1 _10326_/X sky130_fd_sc_hd__mux2_1
X_14094_ _18428_/Q _13834_/X _14092_/X _14093_/X vssd1 vssd1 vccd1 vccd1 _14094_/X
+ sky130_fd_sc_hd__a211o_1
X_18971_ _18972_/CLK _18971_/D vssd1 vssd1 vccd1 vccd1 _18971_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_98_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13045_ _17994_/Q _12783_/A _13025_/A _13041_/Y _11025_/B vssd1 vssd1 vccd1 vccd1
+ _13046_/B sky130_fd_sc_hd__a32o_1
X_17922_ _18988_/CLK _17922_/D vssd1 vssd1 vccd1 vccd1 _17922_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_3_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10257_ _18128_/Q _10257_/B vssd1 vssd1 vccd1 vccd1 _11916_/A sky130_fd_sc_hd__xnor2_1
XFILLER_78_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17853_ _17891_/CLK _17853_/D vssd1 vssd1 vccd1 vccd1 _17853_/Q sky130_fd_sc_hd__dfxtp_1
X_10188_ _10186_/X _10188_/B vssd1 vssd1 vccd1 vccd1 _10189_/B sky130_fd_sc_hd__and2b_1
XFILLER_121_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_208_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16804_ _16803_/B _16802_/X _16803_/Y _16800_/X vssd1 vssd1 vccd1 vccd1 _18770_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_38_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14996_ _14995_/B _14994_/X _14995_/Y _14980_/X vssd1 vssd1 vccd1 vccd1 _18338_/D
+ sky130_fd_sc_hd__o211a_1
X_17784_ _18125_/CLK _17784_/D vssd1 vssd1 vccd1 vccd1 _17784_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_208_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_219_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16735_ _18789_/Q _18753_/Q _16742_/S vssd1 vssd1 vccd1 vccd1 _16735_/X sky130_fd_sc_hd__mux2_1
X_13947_ _18802_/Q _13940_/X _13730_/X _18805_/Q _13946_/X vssd1 vssd1 vccd1 vccd1
+ _13947_/X sky130_fd_sc_hd__a221o_2
XFILLER_47_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_223_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16666_ _16678_/A _16666_/B _16716_/C vssd1 vssd1 vccd1 vccd1 _16666_/X sky130_fd_sc_hd__or3_1
XFILLER_62_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13878_ _18901_/Q _13560_/A _13739_/X _18892_/Q vssd1 vssd1 vccd1 vccd1 _13878_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_228_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15617_ _18484_/Q _15618_/B _15615_/Y _15616_/X vssd1 vssd1 vccd1 vccd1 _18484_/D
+ sky130_fd_sc_hd__o211a_1
X_18405_ _18406_/CLK _18405_/D vssd1 vssd1 vccd1 vccd1 _18405_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_201_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12829_ _17967_/Q vssd1 vssd1 vccd1 vccd1 _12913_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_16597_ _16599_/B _16595_/X _16596_/Y _16581_/X vssd1 vssd1 vccd1 vccd1 _18718_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_98_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15548_ _15993_/A _15548_/B vssd1 vssd1 vccd1 vccd1 _15558_/B sky130_fd_sc_hd__nor2_1
XFILLER_194_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18336_ _18343_/CLK _18336_/D vssd1 vssd1 vccd1 vccd1 _18336_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_1290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_187_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_175_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_1178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18267_ _18275_/CLK _18267_/D vssd1 vssd1 vccd1 vccd1 _18267_/Q sky130_fd_sc_hd__dfxtp_1
X_15479_ _15568_/A vssd1 vssd1 vccd1 vccd1 _15494_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_30_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17218_ _17323_/A vssd1 vssd1 vccd1 vccd1 _17304_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_198_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18198_ _18203_/CLK _18198_/D vssd1 vssd1 vccd1 vccd1 _18198_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_156_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_190_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17149_ _17193_/A _17437_/B _17173_/C vssd1 vssd1 vccd1 vccd1 _17149_/X sky130_fd_sc_hd__or3_1
XFILLER_115_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_196_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09971_ _09386_/A _09376_/B _09971_/S vssd1 vssd1 vccd1 vccd1 _09971_/X sky130_fd_sc_hd__mux2_1
XFILLER_170_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_226_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_1299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_214_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_225_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_1_0_1_wb_clk_i clkbuf_1_0_1_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_2_1_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_168_1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09405_ _18323_/Q _18322_/Q _18321_/Q vssd1 vssd1 vccd1 vccd1 _09408_/B sky130_fd_sc_hd__or3_2
XFILLER_52_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_197_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09336_ _18551_/Q _18550_/Q _18549_/Q vssd1 vssd1 vccd1 vccd1 _09337_/D sky130_fd_sc_hd__or3_4
XFILLER_179_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_221_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09267_ _18965_/Q _18964_/Q _18963_/Q vssd1 vssd1 vccd1 vccd1 _09270_/B sky130_fd_sc_hd__or3_2
XFILLER_166_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09198_ _09198_/A _09198_/B _09198_/C _10293_/A vssd1 vssd1 vccd1 vccd1 _09204_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_5_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11160_ _11160_/A vssd1 vssd1 vccd1 vccd1 _17804_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_84_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10111_ _10032_/X _10068_/X _10109_/X _10110_/Y vssd1 vssd1 vccd1 vccd1 _13410_/C
+ sky130_fd_sc_hd__o31a_1
XFILLER_121_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11091_ _11974_/B _11892_/A _11091_/S vssd1 vssd1 vccd1 vccd1 _11092_/A sky130_fd_sc_hd__mux2_1
XFILLER_175_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10042_ _10086_/A _10035_/X _10037_/X _10069_/A _10076_/S vssd1 vssd1 vccd1 vccd1
+ _10042_/X sky130_fd_sc_hd__a221o_1
XTAP_5534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_216_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_212_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14850_ _14849_/B _14848_/X _14849_/Y _14839_/X vssd1 vssd1 vccd1 vccd1 _18302_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_76_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13801_ _18363_/Q _13670_/X _13743_/A _18339_/Q vssd1 vssd1 vccd1 vccd1 _13801_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_217_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14781_ _18321_/Q _18285_/Q _14787_/S vssd1 vssd1 vccd1 vccd1 _14781_/X sky130_fd_sc_hd__mux2_1
XFILLER_21_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11993_ _14307_/A _13635_/A vssd1 vssd1 vccd1 vccd1 _11993_/X sky130_fd_sc_hd__xor2_2
XFILLER_217_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_216_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16520_ _18699_/Q _16525_/B _16518_/X _16519_/X vssd1 vssd1 vccd1 vccd1 _18699_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_217_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13732_ _13780_/A vssd1 vssd1 vccd1 vccd1 _13732_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_28_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10944_ _09418_/B _09413_/C _10944_/S vssd1 vssd1 vccd1 vccd1 _10944_/X sky130_fd_sc_hd__mux2_1
XFILLER_45_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_231_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_91_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16451_ _16450_/B _16449_/X _16450_/Y _16437_/X vssd1 vssd1 vccd1 vccd1 _18683_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_147_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13663_ _13738_/A vssd1 vssd1 vccd1 vccd1 _13663_/X sky130_fd_sc_hd__buf_8
XFILLER_95_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_1268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10875_ _09392_/C _09397_/B _09402_/D _09397_/D _10695_/X _10856_/S vssd1 vssd1 vccd1
+ vccd1 _10875_/X sky130_fd_sc_hd__mux4_1
XFILLER_71_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_231_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_223_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15402_ _18470_/Q _18434_/Q _15412_/S vssd1 vssd1 vccd1 vccd1 _15402_/X sky130_fd_sc_hd__mux2_1
XFILLER_31_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_227_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_176_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19170_ _19170_/A _09018_/Y vssd1 vssd1 vccd1 vccd1 io_out[8] sky130_fd_sc_hd__ebufn_8
X_12614_ _12609_/B _12523_/X _12613_/Y _12510_/X vssd1 vssd1 vccd1 vccd1 _17925_/D
+ sky130_fd_sc_hd__a211o_1
X_16382_ _16493_/A vssd1 vssd1 vccd1 vccd1 _16473_/A sky130_fd_sc_hd__clkbuf_2
XPHY_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13594_ _13594_/A vssd1 vssd1 vccd1 vccd1 _13705_/A sky130_fd_sc_hd__buf_4
XFILLER_12_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_223_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_85_wb_clk_i _18144_/CLK vssd1 vssd1 vccd1 vccd1 _18593_/CLK sky130_fd_sc_hd__clkbuf_16
XPHY_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18121_ _19028_/CLK _18121_/D vssd1 vssd1 vccd1 vccd1 _18121_/Q sky130_fd_sc_hd__dfxtp_1
X_15333_ _15339_/B _15330_/X _15332_/X _15315_/X vssd1 vssd1 vccd1 vccd1 _18417_/D
+ sky130_fd_sc_hd__o211a_1
XPHY_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12545_ _12556_/A _12542_/Y _12544_/X vssd1 vssd1 vccd1 vccd1 _12545_/X sky130_fd_sc_hd__a21o_1
XFILLER_184_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_185_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_223_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_14_wb_clk_i clkbuf_5_5_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18862_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_18052_ _18052_/CLK _18052_/D vssd1 vssd1 vccd1 vccd1 _18052_/Q sky130_fd_sc_hd__dfxtp_1
X_15264_ _15283_/A vssd1 vssd1 vccd1 vccd1 _15264_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_129_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12476_ _12486_/B _12476_/B vssd1 vssd1 vccd1 vccd1 _12476_/X sky130_fd_sc_hd__and2_1
XFILLER_172_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17003_ _17015_/A _17437_/B _17028_/C vssd1 vssd1 vccd1 vccd1 _17003_/X sky130_fd_sc_hd__or3_1
XFILLER_32_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14215_ _14212_/X _14213_/Y _14214_/Y vssd1 vssd1 vccd1 vccd1 _14342_/B sky130_fd_sc_hd__a21o_1
X_11427_ _11431_/A _17882_/Q _17881_/Q vssd1 vssd1 vccd1 vccd1 _11428_/B sky130_fd_sc_hd__nor3_2
X_15195_ _15239_/A _15195_/B vssd1 vssd1 vccd1 vccd1 _15195_/Y sky130_fd_sc_hd__nand2_1
XFILLER_126_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_193_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14146_ _18560_/Q _14019_/A _13592_/X _18584_/Q vssd1 vssd1 vccd1 vccd1 _14146_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_126_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11358_ _11586_/A vssd1 vssd1 vccd1 vccd1 _11503_/A sky130_fd_sc_hd__inv_2
XFILLER_98_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_193_1277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10309_ _09160_/C _10375_/S _10308_/X _09905_/A vssd1 vssd1 vccd1 vccd1 _10309_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_193_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14077_ _18719_/Q _13596_/X _13630_/X _18701_/Q vssd1 vssd1 vccd1 vccd1 _14077_/X
+ sky130_fd_sc_hd__a22o_1
X_18954_ _18959_/CLK _18954_/D vssd1 vssd1 vccd1 vccd1 _18954_/Q sky130_fd_sc_hd__dfxtp_2
X_11289_ _11286_/X _11617_/A _11661_/A vssd1 vssd1 vccd1 vccd1 _11289_/X sky130_fd_sc_hd__o21a_1
XFILLER_98_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17905_ _17907_/CLK _17905_/D vssd1 vssd1 vccd1 vccd1 _17905_/Q sky130_fd_sc_hd__dfxtp_1
X_13028_ _17987_/Q _13036_/B vssd1 vssd1 vccd1 vccd1 _13028_/X sky130_fd_sc_hd__or2_1
XFILLER_100_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_230_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18885_ _18893_/CLK _18885_/D vssd1 vssd1 vccd1 vccd1 _18885_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_227_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_230_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_227_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17836_ _18209_/CLK _17836_/D vssd1 vssd1 vccd1 vccd1 _17836_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_13_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17767_ _10155_/A _13337_/A _13368_/Y vssd1 vssd1 vccd1 vccd1 _17768_/C sky130_fd_sc_hd__a21o_1
XFILLER_94_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14979_ _14992_/A _14983_/B vssd1 vssd1 vccd1 vccd1 _14979_/Y sky130_fd_sc_hd__nand2_1
XFILLER_19_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16718_ _16766_/A vssd1 vssd1 vccd1 vccd1 _16742_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_207_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_1316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17698_ _17779_/Q _14383_/B _14404_/X vssd1 vssd1 vccd1 vccd1 _17698_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_222_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16649_ _16648_/B _16646_/X _16648_/Y _16639_/X vssd1 vssd1 vccd1 vccd1 _18731_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_222_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_210_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09121_ _09121_/A _09120_/Y vssd1 vssd1 vccd1 vccd1 _09138_/A sky130_fd_sc_hd__or2b_1
XFILLER_194_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18319_ _18324_/CLK _18319_/D vssd1 vssd1 vccd1 vccd1 _18319_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_37_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_202_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09052_ _09052_/A vssd1 vssd1 vccd1 vccd1 _09052_/Y sky130_fd_sc_hd__inv_2
XFILLER_124_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_190_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09954_ _09402_/B _09950_/X _09952_/X _09969_/A vssd1 vssd1 vccd1 vccd1 _09954_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_103_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_132_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_213_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09885_ _09939_/A _09939_/B vssd1 vssd1 vccd1 vccd1 _09974_/A sky130_fd_sc_hd__xor2_4
XFILLER_100_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_213_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_214_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10660_ _10858_/S vssd1 vssd1 vccd1 vccd1 _10660_/X sky130_fd_sc_hd__buf_4
XFILLER_41_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09319_ _09319_/A _09319_/B _09319_/C _09319_/D vssd1 vssd1 vccd1 vccd1 _09320_/C
+ sky130_fd_sc_hd__and4_1
XFILLER_210_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10591_ _09332_/A _09327_/A _09337_/B _10782_/A _10024_/A _10568_/X vssd1 vssd1 vccd1
+ vccd1 _10591_/X sky130_fd_sc_hd__mux4_1
XFILLER_220_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12330_ _12330_/A _12347_/B _12330_/C vssd1 vssd1 vccd1 vccd1 _12331_/A sky130_fd_sc_hd__and3_1
XFILLER_127_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_215_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_193_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12261_ _12261_/A _12261_/B vssd1 vssd1 vccd1 vccd1 _12261_/Y sky130_fd_sc_hd__nor2_1
XFILLER_181_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_218_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14000_ _18937_/Q _13559_/A _13735_/A _18919_/Q vssd1 vssd1 vccd1 vccd1 _14000_/X
+ sky130_fd_sc_hd__a22o_1
X_11212_ _13094_/A _11212_/B vssd1 vssd1 vccd1 vccd1 _11243_/A sky130_fd_sc_hd__nor2_1
XFILLER_134_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12192_ _17897_/Q _17896_/Q _17895_/Q _17894_/Q vssd1 vssd1 vccd1 vccd1 _12193_/D
+ sky130_fd_sc_hd__or4_1
XFILLER_123_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11143_ _11681_/D _17811_/Q _11149_/S vssd1 vssd1 vccd1 vccd1 _11144_/A sky130_fd_sc_hd__mux2_1
XTAP_6021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_6032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_6043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_132_wb_clk_i clkbuf_5_24_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18380_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_66_1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11074_ _17789_/Q vssd1 vssd1 vccd1 vccd1 _11975_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_95_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15951_ _15951_/A vssd1 vssd1 vccd1 vccd1 _17222_/A sky130_fd_sc_hd__buf_8
XTAP_6076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14902_ _14980_/A vssd1 vssd1 vccd1 vccd1 _14902_/X sky130_fd_sc_hd__clkbuf_2
X_10025_ _10025_/A vssd1 vssd1 vccd1 vccd1 _10025_/X sky130_fd_sc_hd__buf_2
XFILLER_209_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18670_ _18686_/CLK _18670_/D vssd1 vssd1 vccd1 vccd1 _18670_/Q sky130_fd_sc_hd__dfxtp_4
XTAP_5364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15882_ _15890_/B _15879_/X _15880_/X _15881_/X vssd1 vssd1 vccd1 vccd1 _18549_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_7_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17621_ _17616_/Y _17561_/X _18968_/Q vssd1 vssd1 vccd1 vccd1 _17621_/X sky130_fd_sc_hd__a21o_1
X_14833_ _14833_/A vssd1 vssd1 vccd1 vccd1 _14848_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_36_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14764_ _14767_/B _14761_/X _14763_/Y _14758_/X vssd1 vssd1 vccd1 vccd1 _18280_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_17_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17552_ _17552_/A vssd1 vssd1 vccd1 vccd1 _17552_/X sky130_fd_sc_hd__clkbuf_2
XTAP_3984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11976_ _11976_/A _11976_/B _12020_/A vssd1 vssd1 vccd1 vccd1 _12025_/D sky130_fd_sc_hd__and3_1
XFILLER_204_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16503_ _16503_/A vssd1 vssd1 vccd1 vccd1 _16555_/A sky130_fd_sc_hd__clkbuf_2
X_13715_ _13715_/A vssd1 vssd1 vccd1 vccd1 _13715_/X sky130_fd_sc_hd__buf_6
X_10927_ _09332_/B _09327_/B _09337_/C _09327_/C _10412_/A _10411_/A vssd1 vssd1 vccd1
+ vccd1 _10927_/X sky130_fd_sc_hd__mux4_1
X_17483_ _17493_/A _17483_/B _17516_/C vssd1 vssd1 vccd1 vccd1 _17483_/X sky130_fd_sc_hd__or3_1
X_14695_ _14944_/A vssd1 vssd1 vccd1 vccd1 _14750_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_60_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_220_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19222_ _19222_/A _08956_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[22] sky130_fd_sc_hd__ebufn_8
XFILLER_108_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16434_ _16434_/A _16880_/B _16481_/C vssd1 vssd1 vccd1 vccd1 _16434_/X sky130_fd_sc_hd__or3_1
XFILLER_147_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13646_ _18885_/Q _14016_/A _13639_/X _13645_/X vssd1 vssd1 vccd1 vccd1 _13646_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_158_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10858_ _09418_/C _09413_/D _10858_/S vssd1 vssd1 vccd1 vccd1 _10858_/X sky130_fd_sc_hd__mux2_1
XFILLER_60_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16365_ _16364_/B _16363_/X _16364_/Y _16354_/X vssd1 vssd1 vccd1 vccd1 _18662_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_176_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19153_ _19153_/A _08954_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[23] sky130_fd_sc_hd__ebufn_8
XFILLER_31_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_160_1243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13577_ _14016_/A vssd1 vssd1 vccd1 vccd1 _13577_/X sky130_fd_sc_hd__buf_2
X_10789_ _09294_/A _09304_/B _10569_/A _09294_/D _10813_/B _10668_/A vssd1 vssd1 vccd1
+ vccd1 _10790_/C sky130_fd_sc_hd__mux4_1
XPHY_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15316_ _15325_/B _15310_/X _15312_/X _15315_/X vssd1 vssd1 vccd1 vccd1 _18414_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_118_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18104_ _18110_/CLK _18104_/D vssd1 vssd1 vccd1 vccd1 _18104_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_185_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12528_ _18132_/Q _15015_/B _12528_/C vssd1 vssd1 vccd1 vccd1 _12591_/A sky130_fd_sc_hd__and3_2
X_16296_ _18644_/Q _16294_/B _16294_/Y _16295_/X vssd1 vssd1 vccd1 vccd1 _18644_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_118_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15247_ _15247_/A vssd1 vssd1 vccd1 vccd1 _15301_/A sky130_fd_sc_hd__buf_2
XFILLER_184_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18035_ _18035_/CLK _18035_/D vssd1 vssd1 vccd1 vccd1 _18035_/Q sky130_fd_sc_hd__dfxtp_1
X_12459_ _12459_/A _12459_/B _12459_/C vssd1 vssd1 vccd1 vccd1 _12460_/A sky130_fd_sc_hd__and3_1
XFILLER_173_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15178_ _15178_/A _15182_/B vssd1 vssd1 vccd1 vccd1 _15178_/Y sky130_fd_sc_hd__nand2_1
XFILLER_99_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14129_ _18290_/Q _13561_/A _13858_/A _18281_/Q vssd1 vssd1 vccd1 vccd1 _14129_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_67_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18937_ _18965_/CLK _18937_/D vssd1 vssd1 vccd1 vccd1 _18937_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_101_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09670_ _09668_/A _09640_/B _09669_/X vssd1 vssd1 vccd1 vccd1 _12070_/B sky130_fd_sc_hd__a21oi_2
XFILLER_28_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18868_ _18870_/CLK _18868_/D vssd1 vssd1 vccd1 vccd1 _18868_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_227_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_223_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_228_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17819_ _17821_/CLK _17819_/D vssd1 vssd1 vccd1 vccd1 _17819_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18799_ _18799_/CLK _18799_/D vssd1 vssd1 vccd1 vccd1 _18799_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_54_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_223_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINSDIODE2_250 _09103_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_261 _14019_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_223_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_272 _18316_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_206_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09104_ _09104_/A _09104_/B _09104_/C vssd1 vssd1 vccd1 vccd1 _09121_/A sky130_fd_sc_hd__and3_1
XFILLER_202_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_182_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19117__88 vssd1 vssd1 vccd1 vccd1 _19117__88/HI _19225_/A sky130_fd_sc_hd__conb_1
X_09035_ _09053_/A vssd1 vssd1 vccd1 vccd1 _09040_/A sky130_fd_sc_hd__buf_12
XFILLER_184_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_131_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_1278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_137_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09937_ _09937_/A vssd1 vssd1 vccd1 vccd1 _09937_/X sky130_fd_sc_hd__buf_4
XFILLER_77_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_213_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_219_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09868_ _18124_/Q _09868_/B vssd1 vssd1 vccd1 vccd1 _09876_/A sky130_fd_sc_hd__xor2_2
XFILLER_100_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_213_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09799_ _09802_/B _09749_/C _09749_/B vssd1 vssd1 vccd1 vccd1 _09808_/A sky130_fd_sc_hd__a21bo_1
XTAP_3247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11830_ _13427_/A _13448_/A _11070_/X vssd1 vssd1 vccd1 vccd1 _11830_/X sky130_fd_sc_hd__a21o_1
XTAP_2524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_227_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_165_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11761_ _11761_/A _11761_/B vssd1 vssd1 vccd1 vccd1 _11763_/B sky130_fd_sc_hd__nand2_1
XTAP_1834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_1295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_159_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13500_ _13500_/A vssd1 vssd1 vccd1 vccd1 _13500_/X sky130_fd_sc_hd__buf_4
XTAP_1856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_5_19_0_wb_clk_i clkbuf_4_9_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18254_/CLK
+ sky130_fd_sc_hd__clkbuf_2
X_10712_ _10805_/B vssd1 vssd1 vccd1 vccd1 _10833_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_14_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14480_ _18215_/Q _14480_/B vssd1 vssd1 vccd1 vccd1 _14481_/A sky130_fd_sc_hd__and2_1
XFILLER_57_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11692_ _17852_/Q _17851_/Q vssd1 vssd1 vccd1 vccd1 _11709_/B sky130_fd_sc_hd__or2_1
XTAP_1889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13431_ _13448_/A _13428_/Y _13430_/X vssd1 vssd1 vccd1 vccd1 _13458_/B sky130_fd_sc_hd__o21ai_2
X_10643_ _10737_/S vssd1 vssd1 vccd1 vccd1 _10644_/A sky130_fd_sc_hd__buf_4
XFILLER_42_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_224_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16150_ _16745_/A _16150_/B vssd1 vssd1 vccd1 vccd1 _16160_/B sky130_fd_sc_hd__nor2_2
XFILLER_158_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13362_ _13362_/A vssd1 vssd1 vccd1 vccd1 _18105_/D sky130_fd_sc_hd__clkbuf_1
X_10574_ _09309_/A _09319_/D _10575_/B vssd1 vssd1 vccd1 vccd1 _10574_/X sky130_fd_sc_hd__mux2_1
X_15101_ _15115_/A _15107_/B vssd1 vssd1 vccd1 vccd1 _15101_/Y sky130_fd_sc_hd__nand2_1
XFILLER_158_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12313_ _17879_/Q _12313_/B vssd1 vssd1 vccd1 vccd1 _12314_/A sky130_fd_sc_hd__and2_1
X_16081_ _16216_/A vssd1 vssd1 vccd1 vccd1 _16132_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_182_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13293_ _18065_/Q _18064_/Q _18067_/Q _18066_/Q vssd1 vssd1 vccd1 vccd1 _13298_/A
+ sky130_fd_sc_hd__or4_1
XFILLER_170_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15032_ _15038_/B _15030_/X _15031_/X _15026_/X vssd1 vssd1 vccd1 vccd1 _18345_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_181_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12244_ _11648_/X _12269_/B _12243_/Y _12219_/X vssd1 vssd1 vccd1 vccd1 _17860_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_218_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12175_ _12180_/A _12175_/B vssd1 vssd1 vccd1 vccd1 _12175_/Y sky130_fd_sc_hd__nor2_1
XFILLER_122_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11126_ _11467_/D vssd1 vssd1 vccd1 vccd1 _11455_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_1_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16983_ _17012_/A vssd1 vssd1 vccd1 vccd1 _17028_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_3_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_231_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18722_ _18722_/CLK _18722_/D vssd1 vssd1 vccd1 vccd1 _18722_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_67_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15934_ _16193_/A vssd1 vssd1 vccd1 vccd1 _15984_/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_5150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11057_ _11336_/B vssd1 vssd1 vccd1 vccd1 _13448_/A sky130_fd_sc_hd__clkbuf_2
XTAP_5161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10008_ _10008_/A vssd1 vssd1 vccd1 vccd1 _10009_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_225_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18653_ _18663_/CLK _18653_/D vssd1 vssd1 vccd1 vccd1 _18653_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_5194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15865_ _15876_/A _15865_/B vssd1 vssd1 vccd1 vccd1 _15865_/Y sky130_fd_sc_hd__nand2_1
XTAP_4460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17604_ _17675_/A vssd1 vssd1 vccd1 vccd1 _17604_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_91_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_1176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14816_ _15255_/A _14841_/B vssd1 vssd1 vccd1 vccd1 _14827_/B sky130_fd_sc_hd__nor2_2
X_18584_ _18590_/CLK _18584_/D vssd1 vssd1 vccd1 vccd1 _18584_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_36_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15796_ _15795_/B _15794_/X _15795_/Y _15783_/X vssd1 vssd1 vccd1 vccd1 _18527_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_3770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_229_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17535_ _17534_/B _17533_/X _17534_/Y _11816_/X vssd1 vssd1 vccd1 vccd1 _18947_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_225_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14747_ _14793_/A _15186_/B _14757_/C vssd1 vssd1 vccd1 vccd1 _14747_/X sky130_fd_sc_hd__or3_1
XFILLER_44_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11959_ _11946_/X _11958_/X _11948_/X vssd1 vssd1 vccd1 vccd1 _11960_/B sky130_fd_sc_hd__a21oi_2
XFILLER_83_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_229_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_225_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14678_ _16949_/A vssd1 vssd1 vccd1 vccd1 _15268_/B sky130_fd_sc_hd__buf_6
XFILLER_33_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17466_ _17469_/B _17463_/X _17465_/Y _17461_/X vssd1 vssd1 vccd1 vccd1 _18928_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_178_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_225_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19205_ _19205_/A _08972_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[5] sky130_fd_sc_hd__ebufn_8
XFILLER_60_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16417_ _16450_/A _16417_/B vssd1 vssd1 vccd1 vccd1 _16417_/Y sky130_fd_sc_hd__nand2_1
X_13629_ _18450_/Q _13591_/X _13625_/X _18456_/Q _13628_/X vssd1 vssd1 vccd1 vccd1
+ _13629_/X sky130_fd_sc_hd__a221o_1
XFILLER_203_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17397_ _17536_/A _17397_/B vssd1 vssd1 vccd1 vccd1 _17408_/B sky130_fd_sc_hd__nor2_2
XFILLER_125_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19136_ _19136_/A _09044_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[6] sky130_fd_sc_hd__ebufn_8
XFILLER_192_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16348_ _16348_/A vssd1 vssd1 vccd1 vccd1 _16363_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_160_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16279_ _16521_/A vssd1 vssd1 vccd1 vccd1 _16325_/A sky130_fd_sc_hd__buf_2
XFILLER_12_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18018_ _18224_/CLK _18018_/D vssd1 vssd1 vccd1 vccd1 _18018_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_218_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09722_ _09594_/X _09722_/B vssd1 vssd1 vccd1 vccd1 _09723_/B sky130_fd_sc_hd__and2b_1
XFILLER_68_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09653_ _09653_/A _09653_/B vssd1 vssd1 vccd1 vccd1 _09654_/B sky130_fd_sc_hd__and2_1
XFILLER_67_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_215_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09584_ _09585_/A _09585_/B _09585_/C vssd1 vssd1 vccd1 vccd1 _09586_/A sky130_fd_sc_hd__o21ai_1
XTAP_1108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_231_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_208_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_169_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_223_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_183_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_1282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_195_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09018_ _09022_/A vssd1 vssd1 vccd1 vccd1 _09018_/Y sky130_fd_sc_hd__inv_2
XFILLER_3_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10290_ _09203_/A _09198_/C _09193_/D _09203_/D _10291_/A _09945_/X vssd1 vssd1 vccd1
+ vccd1 _10290_/X sky130_fd_sc_hd__mux4_2
XFILLER_128_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_120_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_219_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13980_ _18364_/Q _13670_/A _13743_/A _18340_/Q vssd1 vssd1 vccd1 vccd1 _13980_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_4_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_219_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_218_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12931_ _12931_/A vssd1 vssd1 vccd1 vccd1 _12955_/A sky130_fd_sc_hd__clkbuf_2
XTAP_3000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_85_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15650_ _15889_/A vssd1 vssd1 vccd1 vccd1 _15694_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_160_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12862_ _12874_/A vssd1 vssd1 vccd1 vccd1 _12862_/X sky130_fd_sc_hd__buf_6
XTAP_2310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14601_ _16865_/A vssd1 vssd1 vccd1 vccd1 _15199_/B sky130_fd_sc_hd__buf_6
X_11813_ _11867_/A vssd1 vssd1 vccd1 vccd1 _11813_/Y sky130_fd_sc_hd__inv_2
XTAP_3088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15581_ _18512_/Q _18476_/Q _15586_/S vssd1 vssd1 vccd1 vccd1 _15581_/X sky130_fd_sc_hd__mux2_1
XFILLER_160_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12793_ _17958_/Q vssd1 vssd1 vccd1 vccd1 _12793_/Y sky130_fd_sc_hd__inv_2
XTAP_2365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14532_ _14584_/A _15150_/B _14584_/B vssd1 vssd1 vccd1 vccd1 _14532_/X sky130_fd_sc_hd__or3_1
XTAP_1653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17320_ _17370_/A vssd1 vssd1 vccd1 vccd1 _17347_/S sky130_fd_sc_hd__clkbuf_2
X_11744_ _11740_/A _11740_/B _11740_/C vssd1 vssd1 vccd1 vccd1 _11826_/B sky130_fd_sc_hd__a21oi_1
XTAP_1664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17251_ _18911_/Q _18875_/Q _17262_/S vssd1 vssd1 vccd1 vccd1 _17251_/X sky130_fd_sc_hd__mux2_1
X_14463_ _14463_/A _14463_/B vssd1 vssd1 vccd1 vccd1 _14464_/B sky130_fd_sc_hd__nor2_1
XFILLER_109_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11675_ _11653_/B _11848_/B _11673_/X _11674_/X vssd1 vssd1 vccd1 vccd1 _11675_/Y
+ sky130_fd_sc_hd__o31ai_1
XFILLER_230_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16202_ _16202_/A _16202_/B vssd1 vssd1 vccd1 vccd1 _16202_/Y sky130_fd_sc_hd__nand2_1
XFILLER_146_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13414_ _18152_/Q _10990_/X _10982_/X hold3/X vssd1 vssd1 vccd1 vccd1 _18152_/D sky130_fd_sc_hd__a22o_1
XFILLER_174_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10626_ _18122_/Q vssd1 vssd1 vccd1 vccd1 _10640_/A sky130_fd_sc_hd__clkinv_2
X_17182_ _17180_/B _17179_/X _17180_/Y _17181_/X vssd1 vssd1 vccd1 vccd1 _18857_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_139_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14394_ _14391_/Y _14386_/Y _14393_/X _18190_/Q vssd1 vssd1 vccd1 vccd1 _14395_/B
+ sky130_fd_sc_hd__a22o_1
X_16133_ _18608_/Q _16132_/B _16132_/Y _16120_/X vssd1 vssd1 vccd1 vccd1 _18608_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_155_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13345_ _18099_/Q _13344_/X _13342_/X _13339_/X vssd1 vssd1 vccd1 vccd1 _18099_/D
+ sky130_fd_sc_hd__o211a_1
X_10557_ _10549_/A _10556_/X _10443_/A vssd1 vssd1 vccd1 vccd1 _10557_/X sky130_fd_sc_hd__o21a_1
XFILLER_154_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16064_ _16064_/A _16064_/B vssd1 vssd1 vccd1 vccd1 _16064_/Y sky130_fd_sc_hd__nand2_1
XFILLER_154_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13276_ _19018_/Q _19017_/Q _19020_/Q _19019_/Q vssd1 vssd1 vccd1 vccd1 _13278_/C
+ sky130_fd_sc_hd__or4_1
XFILLER_6_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10488_ _09153_/D _09148_/D _09143_/C _09148_/B _12032_/A _10454_/X vssd1 vssd1 vccd1
+ vccd1 _10488_/X sky130_fd_sc_hd__mux4_2
X_15015_ _18148_/Q _15015_/B vssd1 vssd1 vccd1 vccd1 _15125_/A sky130_fd_sc_hd__nand2_2
XFILLER_154_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12227_ _12940_/A vssd1 vssd1 vccd1 vccd1 _12517_/A sky130_fd_sc_hd__buf_6
XFILLER_155_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12158_ _12158_/A _12158_/B vssd1 vssd1 vccd1 vccd1 _12158_/X sky130_fd_sc_hd__or2_1
XFILLER_64_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_4_12_0_wb_clk_i clkbuf_3_6_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_5_25_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_151_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11109_ _11359_/B vssd1 vssd1 vccd1 vccd1 _11404_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_110_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16966_ _18841_/Q _18805_/Q _16970_/S vssd1 vssd1 vccd1 vccd1 _16966_/X sky130_fd_sc_hd__mux2_1
X_12089_ _12089_/A _12089_/B vssd1 vssd1 vccd1 vccd1 _12095_/A sky130_fd_sc_hd__xnor2_1
XFILLER_49_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18705_ _18708_/CLK _18705_/D vssd1 vssd1 vccd1 vccd1 _18705_/Q sky130_fd_sc_hd__dfxtp_2
X_15917_ _18142_/Q _16528_/B vssd1 vssd1 vccd1 vccd1 _16034_/A sky130_fd_sc_hd__nand2_2
XFILLER_204_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16897_ _17164_/A vssd1 vssd1 vccd1 vccd1 _16954_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_225_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_37_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18636_ _18641_/CLK _18636_/D vssd1 vssd1 vccd1 vccd1 _18636_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_94_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15848_ _15853_/B _15846_/X _15847_/X _15842_/X vssd1 vssd1 vccd1 vccd1 _18540_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_4290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18567_ _18571_/CLK _18567_/D vssd1 vssd1 vccd1 vccd1 _18567_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_24_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15779_ _15815_/A _15782_/B vssd1 vssd1 vccd1 vccd1 _15779_/Y sky130_fd_sc_hd__nand2_1
XFILLER_212_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_205_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_221_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_178_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17518_ _17524_/B _17515_/X _17516_/X _17517_/X vssd1 vssd1 vccd1 vccd1 _18942_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_127_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18498_ _18504_/CLK _18498_/D vssd1 vssd1 vccd1 vccd1 _18498_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_205_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_221_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17449_ _17493_/A _17449_/B _17460_/C vssd1 vssd1 vccd1 vccd1 _17449_/X sky130_fd_sc_hd__or3_1
XFILLER_220_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_221_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_229_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_229_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_5 _09058_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_214_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09705_ _10568_/A vssd1 vssd1 vccd1 vccd1 _10060_/A sky130_fd_sc_hd__buf_2
XFILLER_74_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_216_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_210_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09636_ _09637_/A _09637_/B vssd1 vssd1 vccd1 vccd1 _09642_/B sky130_fd_sc_hd__xnor2_1
XFILLER_215_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_216_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09567_ _09568_/A _09576_/B vssd1 vssd1 vccd1 vccd1 _09573_/A sky130_fd_sc_hd__xor2_1
XFILLER_231_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_224_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_196_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_230_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09498_ _18196_/Q _09498_/B vssd1 vssd1 vccd1 vccd1 _09499_/B sky130_fd_sc_hd__or2_1
XFILLER_90_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_212_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11460_ _17887_/Q vssd1 vssd1 vccd1 vccd1 _11478_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_7_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10411_ _10411_/A vssd1 vssd1 vccd1 vccd1 _10496_/A sky130_fd_sc_hd__buf_4
XFILLER_104_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_221_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11391_ _11619_/A _11386_/X _11388_/Y _11390_/X vssd1 vssd1 vccd1 vccd1 _11391_/Y
+ sky130_fd_sc_hd__o22ai_1
XFILLER_164_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13130_ _13130_/A vssd1 vssd1 vccd1 vccd1 _18024_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_87_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10342_ _10338_/X _10341_/X _09889_/X vssd1 vssd1 vccd1 vccd1 _10342_/X sky130_fd_sc_hd__o21a_1
XFILLER_99_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13061_ _13375_/B _12776_/X _13060_/Y _13037_/X vssd1 vssd1 vccd1 vccd1 _17997_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_140_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10273_ _09209_/A _09214_/D _10285_/S vssd1 vssd1 vccd1 vccd1 _10273_/X sky130_fd_sc_hd__mux2_1
XFILLER_133_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12012_ _14289_/A _12129_/A vssd1 vssd1 vccd1 vccd1 _12012_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_105_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19101__72 vssd1 vssd1 vccd1 vccd1 _19101__72/HI _19209_/A sky130_fd_sc_hd__conb_1
Xclkbuf_leaf_39_wb_clk_i _18254_/CLK vssd1 vssd1 vccd1 vccd1 _18773_/CLK sky130_fd_sc_hd__clkbuf_16
X_16820_ _16952_/A vssd1 vssd1 vccd1 vccd1 _16928_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_94_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16751_ _18793_/Q _18757_/Q _16762_/S vssd1 vssd1 vccd1 vccd1 _16751_/X sky130_fd_sc_hd__mux2_1
X_13963_ _18433_/Q _13847_/A _13781_/X _18424_/Q vssd1 vssd1 vccd1 vccd1 _13963_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_19_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_219_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15702_ _18541_/Q _18505_/Q _15714_/S vssd1 vssd1 vccd1 vccd1 _15702_/X sky130_fd_sc_hd__mux2_1
XFILLER_111_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12914_ _17966_/Q _12913_/A _12908_/B _17968_/Q vssd1 vssd1 vccd1 vccd1 _12915_/C
+ sky130_fd_sc_hd__a31o_1
XFILLER_185_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13894_ _18610_/Q _13594_/A _13535_/A _18592_/Q vssd1 vssd1 vccd1 vccd1 _13894_/X
+ sky130_fd_sc_hd__a22o_1
X_16682_ _16780_/A vssd1 vssd1 vccd1 vccd1 _16760_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_46_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18421_ _18423_/CLK _18421_/D vssd1 vssd1 vccd1 vccd1 _18421_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_34_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15633_ _15633_/A _15633_/B vssd1 vssd1 vccd1 vccd1 _15633_/Y sky130_fd_sc_hd__nand2_1
XFILLER_46_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12845_ _17945_/Q _17946_/Q _17947_/Q vssd1 vssd1 vccd1 vccd1 _12851_/B sky130_fd_sc_hd__and3_1
XTAP_2140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18352_ _18356_/CLK _18352_/D vssd1 vssd1 vccd1 vccd1 _18352_/Q sky130_fd_sc_hd__dfxtp_4
XTAP_2184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15564_ _15570_/B _15561_/X _15563_/X _15555_/X vssd1 vssd1 vccd1 vccd1 _18471_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_1450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12776_ _12786_/B vssd1 vssd1 vccd1 vccd1 _12776_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17303_ _17336_/A _17303_/B vssd1 vssd1 vccd1 vccd1 _17303_/Y sky130_fd_sc_hd__nand2_1
X_11727_ _11727_/A _17913_/Q vssd1 vssd1 vccd1 vccd1 _11727_/Y sky130_fd_sc_hd__nand2_1
X_14515_ _18229_/Q _14515_/B _14515_/C vssd1 vssd1 vccd1 vccd1 _14515_/Y sky130_fd_sc_hd__nor3_1
X_15495_ _15508_/A _15500_/B vssd1 vssd1 vccd1 vccd1 _15495_/Y sky130_fd_sc_hd__nand2_1
X_18283_ _18290_/CLK _18283_/D vssd1 vssd1 vccd1 vccd1 _18283_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_202_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17234_ _17256_/A _17516_/B _17234_/C vssd1 vssd1 vccd1 vccd1 _17234_/X sky130_fd_sc_hd__or3_1
X_11658_ _11658_/A vssd1 vssd1 vccd1 vccd1 _11659_/D sky130_fd_sc_hd__inv_2
X_14446_ _14404_/A _14445_/B _14423_/A vssd1 vssd1 vccd1 vccd1 _14446_/X sky130_fd_sc_hd__a21o_1
XFILLER_168_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10609_ _10731_/A vssd1 vssd1 vccd1 vccd1 _10616_/A sky130_fd_sc_hd__inv_2
XFILLER_127_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14377_ _14377_/A vssd1 vssd1 vccd1 vccd1 _17766_/A sky130_fd_sc_hd__buf_6
X_17165_ _17210_/A _17169_/B vssd1 vssd1 vccd1 vccd1 _17165_/Y sky130_fd_sc_hd__nand2_1
X_11589_ _11297_/B _11588_/X _11313_/B vssd1 vssd1 vccd1 vccd1 _11592_/C sky130_fd_sc_hd__a21oi_1
XFILLER_143_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16116_ _16123_/B _16113_/X _16115_/X _16097_/X vssd1 vssd1 vccd1 vccd1 _18603_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_183_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13328_ _18093_/Q _13313_/X _13327_/Y _13074_/X vssd1 vssd1 vccd1 vccd1 _18093_/D
+ sky130_fd_sc_hd__o211a_1
Xclkbuf_2_2_1_wb_clk_i clkbuf_2_2_1_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_5_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_2
X_17096_ _17096_/A vssd1 vssd1 vccd1 vccd1 _17096_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_192_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16047_ _16273_/A vssd1 vssd1 vccd1 vccd1 _16139_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_171_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13259_ _13259_/A vssd1 vssd1 vccd1 vccd1 _18082_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_171_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_229_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_229_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17998_ _18997_/CLK _17998_/D vssd1 vssd1 vccd1 vccd1 _17998_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16949_ _16949_/A vssd1 vssd1 vccd1 vccd1 _17528_/B sky130_fd_sc_hd__buf_4
Xclkbuf_5_1_0_wb_clk_i clkbuf_5_1_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _17929_/CLK
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_92_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09421_ _09421_/A vssd1 vssd1 vccd1 vccd1 _09421_/Y sky130_fd_sc_hd__inv_2
XFILLER_53_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18619_ _18620_/CLK _18619_/D vssd1 vssd1 vccd1 vccd1 _18619_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_213_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09352_ _18416_/Q _18415_/Q _18414_/Q vssd1 vssd1 vccd1 vccd1 _09354_/C sky130_fd_sc_hd__or3_4
XFILLER_80_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09283_ _18857_/Q _18856_/Q _18855_/Q vssd1 vssd1 vccd1 vccd1 _09287_/A sky130_fd_sc_hd__or3_4
XFILLER_178_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_221_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_173_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_173_1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08998_ _08998_/A vssd1 vssd1 vccd1 vccd1 _09003_/A sky130_fd_sc_hd__buf_12
XTAP_5749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10960_ _09360_/A _09370_/A _09365_/C _09360_/B _09683_/X _09709_/X vssd1 vssd1 vccd1
+ vccd1 _10960_/X sky130_fd_sc_hd__mux4_2
XFILLER_18_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_216_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09619_ _09664_/A vssd1 vssd1 vccd1 vccd1 _09684_/A sky130_fd_sc_hd__buf_2
X_10891_ _09376_/A _09386_/B _09381_/A _09376_/D _10103_/B _10025_/A vssd1 vssd1 vccd1
+ vccd1 _10891_/X sky130_fd_sc_hd__mux4_1
XFILLER_203_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_216_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12630_ _17929_/Q _12630_/B vssd1 vssd1 vccd1 vccd1 _12630_/X sky130_fd_sc_hd__or2_1
XFILLER_31_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_180_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12561_ _17923_/Q _12570_/B vssd1 vssd1 vccd1 vccd1 _12561_/Y sky130_fd_sc_hd__nand2_2
XFILLER_54_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11512_ _19031_/Q _17873_/Q _11512_/C vssd1 vssd1 vccd1 vccd1 _11534_/A sky130_fd_sc_hd__and3_1
X_14300_ _14300_/A vssd1 vssd1 vccd1 vccd1 _14300_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_15280_ _15286_/B _15278_/X _15279_/X _15264_/X vssd1 vssd1 vccd1 vccd1 _18408_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_211_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12492_ _12492_/A vssd1 vssd1 vccd1 vccd1 _12495_/B sky130_fd_sc_hd__inv_2
XFILLER_200_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14231_ _13409_/X _14227_/X _14229_/X _17709_/B _18169_/Q vssd1 vssd1 vccd1 vccd1
+ _14231_/X sky130_fd_sc_hd__a311o_1
XFILLER_172_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11443_ _11795_/A _11788_/A _11732_/A _11652_/B vssd1 vssd1 vccd1 vccd1 _11443_/X
+ sky130_fd_sc_hd__and4_1
XFILLER_109_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14162_ _18956_/Q _14019_/X _13582_/X _18962_/Q vssd1 vssd1 vccd1 vccd1 _14162_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_152_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11374_ _11374_/A _11374_/B _11374_/C vssd1 vssd1 vccd1 vccd1 _11374_/X sky130_fd_sc_hd__and3_1
XFILLER_152_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13113_ _13113_/A vssd1 vssd1 vccd1 vccd1 _18016_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_30_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10325_ _09253_/A _09248_/C _09243_/D _09253_/D _10291_/A _09971_/S vssd1 vssd1 vccd1
+ vccd1 _10325_/X sky130_fd_sc_hd__mux4_1
X_14093_ _18443_/Q _13617_/A _13732_/X _18437_/Q vssd1 vssd1 vccd1 vccd1 _14093_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_152_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18970_ _18970_/CLK _18970_/D vssd1 vssd1 vccd1 vccd1 _18970_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_106_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19078__49 vssd1 vssd1 vccd1 vccd1 _19078__49/HI _19172_/A sky130_fd_sc_hd__conb_1
XFILLER_112_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13044_ _13044_/A vssd1 vssd1 vccd1 vccd1 _17993_/D sky130_fd_sc_hd__clkbuf_1
X_17921_ _17926_/CLK _17921_/D vssd1 vssd1 vccd1 vccd1 _17921_/Q sky130_fd_sc_hd__dfxtp_1
X_10256_ _10256_/A _11913_/S vssd1 vssd1 vccd1 vccd1 _10257_/B sky130_fd_sc_hd__xnor2_1
XFILLER_133_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17852_ _17891_/CLK _17852_/D vssd1 vssd1 vccd1 vccd1 _17852_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_66_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10187_ _18100_/Q _10623_/A vssd1 vssd1 vccd1 vccd1 _10188_/B sky130_fd_sc_hd__or2_1
XFILLER_117_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16803_ _16815_/A _16803_/B vssd1 vssd1 vccd1 vccd1 _16803_/Y sky130_fd_sc_hd__nand2_1
XFILLER_78_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17783_ _19028_/CLK _17783_/D vssd1 vssd1 vccd1 vccd1 _17783_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_208_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14995_ _14995_/A _14995_/B vssd1 vssd1 vccd1 vccd1 _14995_/Y sky130_fd_sc_hd__nand2_1
XFILLER_94_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16734_ _16734_/A _16745_/B vssd1 vssd1 vccd1 vccd1 _16743_/B sky130_fd_sc_hd__nor2_2
XFILLER_35_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13946_ _18778_/Q _13749_/X _13942_/X _13945_/X vssd1 vssd1 vccd1 vccd1 _13946_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_228_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16665_ _16794_/B vssd1 vssd1 vccd1 vccd1 _16716_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_13877_ _13877_/A vssd1 vssd1 vccd1 vccd1 _13877_/X sky130_fd_sc_hd__buf_12
XFILLER_46_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_223_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18404_ _18404_/CLK _18404_/D vssd1 vssd1 vccd1 vccd1 _18404_/Q sky130_fd_sc_hd__dfxtp_2
X_15616_ _15616_/A vssd1 vssd1 vccd1 vccd1 _15616_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_50_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_222_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12828_ _12588_/B _17951_/Q _17952_/Q _12594_/B _12827_/Y vssd1 vssd1 vccd1 vccd1
+ _12835_/B sky130_fd_sc_hd__o221ai_1
X_16596_ _16631_/A _16599_/B vssd1 vssd1 vccd1 vccd1 _16596_/Y sky130_fd_sc_hd__nand2_1
XFILLER_201_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18335_ _18373_/CLK _18335_/D vssd1 vssd1 vccd1 vccd1 _18335_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_72_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_231_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15547_ _15546_/B _15545_/X _15546_/Y _15536_/X vssd1 vssd1 vccd1 vccd1 _18467_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_1280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12759_ _12919_/B _12921_/B _12920_/A _12757_/X _12758_/X vssd1 vssd1 vccd1 vccd1
+ _13318_/B sky130_fd_sc_hd__a41o_2
XTAP_1291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_1277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18266_ _18266_/CLK _18266_/D vssd1 vssd1 vccd1 vccd1 _18266_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_198_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15478_ _15589_/A vssd1 vssd1 vccd1 vccd1 _15568_/A sky130_fd_sc_hd__buf_2
XFILLER_129_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17217_ _17256_/A _17506_/B _17234_/C vssd1 vssd1 vccd1 vccd1 _17217_/X sky130_fd_sc_hd__or3_1
X_14429_ _18197_/Q _14427_/X _14428_/X _09500_/B vssd1 vssd1 vccd1 vccd1 _14430_/B
+ sky130_fd_sc_hd__o2bb2a_1
X_18197_ _18203_/CLK _18197_/D vssd1 vssd1 vccd1 vccd1 _18197_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_128_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17148_ _17148_/A vssd1 vssd1 vccd1 vccd1 _17193_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_196_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09970_ _10292_/S vssd1 vssd1 vccd1 vccd1 _09971_/S sky130_fd_sc_hd__buf_4
XFILLER_116_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17079_ _18869_/Q _18833_/Q _17094_/S vssd1 vssd1 vccd1 vccd1 _17079_/X sky130_fd_sc_hd__mux2_1
XFILLER_171_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_226_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19092__63 vssd1 vssd1 vccd1 vccd1 _19092__63/HI _19200_/A sky130_fd_sc_hd__conb_1
XFILLER_211_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_214_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09404_ _18329_/Q _18328_/Q _18327_/Q vssd1 vssd1 vccd1 vccd1 _09408_/A sky130_fd_sc_hd__or3_2
XFILLER_52_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_213_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_197_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_209_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09335_ _18542_/Q _18541_/Q _18540_/Q vssd1 vssd1 vccd1 vccd1 _09337_/C sky130_fd_sc_hd__or3_2
XFILLER_40_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_1355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_178_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_205_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09266_ _18974_/Q _18973_/Q _18972_/Q vssd1 vssd1 vccd1 vccd1 _09270_/A sky130_fd_sc_hd__or3_2
XFILLER_142_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09197_ _18557_/Q _18556_/Q _18555_/Q vssd1 vssd1 vccd1 vccd1 _10293_/A sky130_fd_sc_hd__or3_4
XFILLER_101_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10110_ _10110_/A vssd1 vssd1 vccd1 vccd1 _10110_/Y sky130_fd_sc_hd__inv_2
XFILLER_171_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11090_ _11963_/A vssd1 vssd1 vccd1 vccd1 _11974_/B sky130_fd_sc_hd__clkbuf_2
XTAP_5502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_1326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10041_ _10041_/A vssd1 vssd1 vccd1 vccd1 _10076_/S sky130_fd_sc_hd__buf_4
XTAP_5524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_216_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_195_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13800_ _18342_/Q _13719_/A _13752_/A _18348_/Q vssd1 vssd1 vccd1 vccd1 _13800_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_4878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14780_ _15218_/A _14790_/B vssd1 vssd1 vccd1 vccd1 _14788_/B sky130_fd_sc_hd__nor2_1
XFILLER_17_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11992_ _12102_/B vssd1 vssd1 vccd1 vccd1 _13635_/A sky130_fd_sc_hd__buf_2
XFILLER_90_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_217_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13731_ _13731_/A vssd1 vssd1 vccd1 vccd1 _13780_/A sky130_fd_sc_hd__clkbuf_4
X_10943_ _09402_/D _10069_/X _10940_/X _09370_/C _10948_/S vssd1 vssd1 vccd1 vccd1
+ _10943_/X sky130_fd_sc_hd__a221o_1
XFILLER_21_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_217_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16450_ _16450_/A _16450_/B vssd1 vssd1 vccd1 vccd1 _16450_/Y sky130_fd_sc_hd__nand2_1
X_10874_ _10757_/A _10869_/X _10873_/X _10733_/X vssd1 vssd1 vccd1 vccd1 _10874_/X
+ sky130_fd_sc_hd__o211a_1
X_13662_ _18984_/Q _14081_/B _13532_/A _18975_/Q _13661_/X vssd1 vssd1 vccd1 vccd1
+ _13662_/X sky130_fd_sc_hd__a221o_1
XFILLER_44_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15401_ _15403_/B _15399_/X _15400_/Y _15382_/X vssd1 vssd1 vccd1 vccd1 _18433_/D
+ sky130_fd_sc_hd__o211a_1
XPHY_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12613_ _12613_/A _12613_/B vssd1 vssd1 vccd1 vccd1 _12613_/Y sky130_fd_sc_hd__nor2_1
XFILLER_231_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_223_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13593_ _18702_/Q _13591_/X _13592_/X _18726_/Q vssd1 vssd1 vccd1 vccd1 _13593_/X
+ sky130_fd_sc_hd__a22o_1
XPHY_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16381_ _18139_/Q _16528_/B vssd1 vssd1 vccd1 vccd1 _16493_/A sky130_fd_sc_hd__nand2_2
XFILLER_31_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18120_ _18130_/CLK _18120_/D vssd1 vssd1 vccd1 vccd1 _18120_/Q sky130_fd_sc_hd__dfxtp_2
X_15332_ _15358_/A _15935_/B _15358_/C vssd1 vssd1 vccd1 vccd1 _15332_/X sky130_fd_sc_hd__or3_1
X_12544_ _12535_/A _12535_/B _12543_/X vssd1 vssd1 vccd1 vccd1 _12544_/X sky130_fd_sc_hd__a21o_1
XFILLER_223_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18051_ _18052_/CLK _18051_/D vssd1 vssd1 vccd1 vccd1 _18051_/Q sky130_fd_sc_hd__dfxtp_1
X_15263_ _15303_/A _15263_/B vssd1 vssd1 vccd1 vccd1 _15263_/Y sky130_fd_sc_hd__nand2_1
X_12475_ _12475_/A vssd1 vssd1 vccd1 vccd1 _12475_/Y sky130_fd_sc_hd__inv_2
XFILLER_184_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17002_ _18849_/Q _18813_/Q _17005_/S vssd1 vssd1 vccd1 vccd1 _17002_/X sky130_fd_sc_hd__mux2_1
XFILLER_8_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11426_ _19029_/Q vssd1 vssd1 vccd1 vccd1 _11431_/A sky130_fd_sc_hd__inv_2
X_14214_ _18211_/Q vssd1 vssd1 vccd1 vccd1 _14214_/Y sky130_fd_sc_hd__inv_2
X_15194_ _15252_/A vssd1 vssd1 vccd1 vccd1 _15239_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_32_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_1204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_54_wb_clk_i _18759_/CLK vssd1 vssd1 vccd1 vccd1 _18752_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_99_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14145_ _18572_/Q _13834_/A _13582_/X _18566_/Q _14144_/X vssd1 vssd1 vccd1 vccd1
+ _14145_/X sky130_fd_sc_hd__a221o_1
X_11357_ _11404_/A _11357_/B vssd1 vssd1 vccd1 vccd1 _11617_/B sky130_fd_sc_hd__nor2_1
XFILLER_67_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10308_ _10308_/A _10376_/B vssd1 vssd1 vccd1 vccd1 _10308_/X sky130_fd_sc_hd__or2_1
XFILLER_3_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14076_ _18704_/Q _13508_/A _13861_/X _18728_/Q vssd1 vssd1 vccd1 vccd1 _14076_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_154_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18953_ _18953_/CLK _18953_/D vssd1 vssd1 vccd1 vccd1 _18953_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_193_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11288_ _11541_/B vssd1 vssd1 vccd1 vccd1 _11617_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_3_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17904_ _17907_/CLK _17904_/D vssd1 vssd1 vccd1 vccd1 _17904_/Q sky130_fd_sc_hd__dfxtp_1
X_13027_ _12975_/A _13025_/X _13026_/X _13011_/X vssd1 vssd1 vccd1 vccd1 _17986_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_112_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10239_ _10466_/A vssd1 vssd1 vccd1 vccd1 _10549_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_67_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18884_ _18907_/CLK _18884_/D vssd1 vssd1 vccd1 vccd1 _18884_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_230_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17835_ _18163_/CLK _17835_/D vssd1 vssd1 vccd1 vccd1 _17835_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_120_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17766_ _17766_/A input6/X vssd1 vssd1 vccd1 vccd1 _19026_/D sky130_fd_sc_hd__nor2_1
X_14978_ _18370_/Q _18334_/Q _14994_/S vssd1 vssd1 vccd1 vccd1 _14978_/X sky130_fd_sc_hd__mux2_1
XFILLER_130_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16717_ _16723_/B _16715_/X _16716_/X _16704_/X vssd1 vssd1 vccd1 vccd1 _18747_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_35_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13929_ _18262_/Q _13615_/A _13927_/X _13928_/X vssd1 vssd1 vccd1 vccd1 _13929_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_78_1355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17697_ _17697_/A vssd1 vssd1 vccd1 vccd1 _18986_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_39_1328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_1208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_222_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16648_ _16699_/A _16648_/B vssd1 vssd1 vccd1 vccd1 _16648_/Y sky130_fd_sc_hd__nand2_1
XFILLER_62_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_222_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16579_ _16615_/A _16880_/B _16628_/C vssd1 vssd1 vccd1 vccd1 _16579_/X sky130_fd_sc_hd__or3_1
XFILLER_176_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09120_ _09120_/A _09120_/B _09120_/C vssd1 vssd1 vccd1 vccd1 _09120_/Y sky130_fd_sc_hd__nand3_1
XFILLER_148_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18318_ _18324_/CLK _18318_/D vssd1 vssd1 vccd1 vccd1 _18318_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_124_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_187_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09051_ _09052_/A vssd1 vssd1 vccd1 vccd1 _09051_/Y sky130_fd_sc_hd__inv_2
XFILLER_191_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18249_ _18251_/CLK _18249_/D vssd1 vssd1 vccd1 vccd1 _18249_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_198_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_191_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_191_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09953_ _09953_/A vssd1 vssd1 vccd1 vccd1 _09969_/A sky130_fd_sc_hd__buf_4
XFILLER_103_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09884_ _09902_/A _09887_/B _09883_/X vssd1 vssd1 vccd1 vccd1 _09939_/B sky130_fd_sc_hd__a21o_4
XFILLER_213_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_213_1348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_218_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09318_ _18461_/Q _18460_/Q _18459_/Q vssd1 vssd1 vccd1 vccd1 _09319_/D sky130_fd_sc_hd__or3_4
XFILLER_167_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10590_ _09337_/A _09332_/C _09327_/D _09337_/D _10046_/A _10568_/X vssd1 vssd1 vccd1
+ vccd1 _10590_/X sky130_fd_sc_hd__mux4_1
XFILLER_16_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09249_ _18890_/Q _18889_/Q _18888_/Q vssd1 vssd1 vccd1 vccd1 _09253_/A sky130_fd_sc_hd__or3_4
XFILLER_31_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12260_ _11563_/B _11556_/X _17869_/Q vssd1 vssd1 vccd1 vccd1 _12261_/B sky130_fd_sc_hd__a21o_1
XFILLER_154_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11211_ _11211_/A vssd1 vssd1 vccd1 vccd1 _17814_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_135_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12191_ _17891_/Q vssd1 vssd1 vccd1 vccd1 _12352_/B sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_6000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11142_ _11795_/A vssd1 vssd1 vccd1 vccd1 _11681_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_218_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19048__19 vssd1 vssd1 vccd1 vccd1 _19048__19/HI _19142_/A sky130_fd_sc_hd__conb_1
XFILLER_123_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_6022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_6033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15950_ _18601_/Q _18565_/Q _15963_/S vssd1 vssd1 vccd1 vccd1 _15950_/X sky130_fd_sc_hd__mux2_1
XTAP_5310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11073_ _11073_/A vssd1 vssd1 vccd1 vccd1 _17788_/D sky130_fd_sc_hd__clkbuf_1
XTAP_5321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14901_ _15207_/A vssd1 vssd1 vccd1 vccd1 _14980_/A sky130_fd_sc_hd__clkbuf_2
X_10024_ _10024_/A vssd1 vssd1 vccd1 vccd1 _10025_/A sky130_fd_sc_hd__buf_4
XTAP_5354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15881_ _15925_/A vssd1 vssd1 vccd1 vccd1 _15881_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_4620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17620_ _14357_/X _14612_/X _17547_/X _17619_/X _17556_/X vssd1 vssd1 vccd1 vccd1
+ _18967_/D sky130_fd_sc_hd__o311a_1
XTAP_5398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14832_ _14838_/B _14830_/X _14831_/X _14819_/X vssd1 vssd1 vccd1 vccd1 _18297_/D
+ sky130_fd_sc_hd__o211a_1
Xclkbuf_leaf_172_wb_clk_i _18114_/CLK vssd1 vssd1 vccd1 vccd1 _18151_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_64_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_101_wb_clk_i clkbuf_5_28_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18548_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_4697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17551_ _17675_/A vssd1 vssd1 vccd1 vccd1 _17552_/A sky130_fd_sc_hd__buf_2
XTAP_3963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14763_ _14810_/A _14767_/B vssd1 vssd1 vccd1 vccd1 _14763_/Y sky130_fd_sc_hd__nand2_1
XFILLER_63_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11975_ _11975_/A _11970_/C vssd1 vssd1 vccd1 vccd1 _12020_/A sky130_fd_sc_hd__or2b_1
XTAP_3985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16502_ _18732_/Q _18696_/Q _16509_/S vssd1 vssd1 vccd1 vccd1 _16502_/X sky130_fd_sc_hd__mux2_1
XTAP_3996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13714_ _13730_/A vssd1 vssd1 vccd1 vccd1 _13714_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_229_1366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17482_ _18969_/Q _18933_/Q _17495_/S vssd1 vssd1 vccd1 vccd1 _17482_/X sky130_fd_sc_hd__mux2_1
X_10926_ _10926_/A _10926_/B vssd1 vssd1 vccd1 vccd1 _10926_/X sky130_fd_sc_hd__and2_1
XFILLER_186_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14694_ _15643_/A vssd1 vssd1 vccd1 vccd1 _14944_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_71_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19221_ _19221_/A _08958_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[21] sky130_fd_sc_hd__ebufn_8
XFILLER_205_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16433_ _16433_/A vssd1 vssd1 vccd1 vccd1 _16481_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_204_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10857_ _09418_/A _09408_/D _10870_/S vssd1 vssd1 vccd1 vccd1 _10857_/X sky130_fd_sc_hd__mux2_1
X_13645_ _18909_/Q _13616_/A _13643_/X _13644_/X vssd1 vssd1 vccd1 vccd1 _13645_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_147_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19152_ _19152_/A _08953_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[22] sky130_fd_sc_hd__ebufn_8
XFILLER_201_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_201_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16364_ _16392_/A _16364_/B vssd1 vssd1 vccd1 vccd1 _16364_/Y sky130_fd_sc_hd__nand2_1
XFILLER_158_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13576_ _13576_/A vssd1 vssd1 vccd1 vccd1 _13576_/X sky130_fd_sc_hd__buf_2
X_10788_ _09337_/A _09332_/C _09327_/D _09337_/D _10701_/A _10883_/B vssd1 vssd1 vccd1
+ vccd1 _10788_/X sky130_fd_sc_hd__mux4_1
XFILLER_9_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_160_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18103_ _18125_/CLK _18103_/D vssd1 vssd1 vccd1 vccd1 _18103_/Q sky130_fd_sc_hd__dfxtp_2
X_15315_ _15404_/A vssd1 vssd1 vccd1 vccd1 _15315_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_157_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12527_ _16673_/A vssd1 vssd1 vccd1 vccd1 _15015_/B sky130_fd_sc_hd__buf_8
X_16295_ _16354_/A vssd1 vssd1 vccd1 vccd1 _16295_/X sky130_fd_sc_hd__clkbuf_2
X_18034_ _18035_/CLK _18034_/D vssd1 vssd1 vccd1 vccd1 _18034_/Q sky130_fd_sc_hd__dfxtp_1
X_15246_ _18436_/Q _18400_/Q _15246_/S vssd1 vssd1 vccd1 vccd1 _15246_/X sky130_fd_sc_hd__mux2_1
XFILLER_173_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_145_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12458_ _12458_/A _12477_/A _12477_/B vssd1 vssd1 vccd1 vccd1 _12459_/C sky130_fd_sc_hd__nand3_1
XFILLER_126_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11409_ _11617_/C _11609_/A vssd1 vssd1 vccd1 vccd1 _11546_/B sky130_fd_sc_hd__nand2_1
X_15177_ _18418_/Q _18382_/Q _15177_/S vssd1 vssd1 vccd1 vccd1 _15177_/X sky130_fd_sc_hd__mux2_1
X_12389_ _12397_/B _12490_/A _12389_/C vssd1 vssd1 vccd1 vccd1 _12390_/A sky130_fd_sc_hd__and3b_1
XFILLER_67_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_154_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14128_ _18914_/Q _14015_/X _14027_/X _18905_/Q _14127_/X vssd1 vssd1 vccd1 vccd1
+ _14128_/X sky130_fd_sc_hd__a221o_1
XFILLER_207_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_1340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14059_ _18398_/Q _13562_/A _13493_/A _18389_/Q _14058_/X vssd1 vssd1 vccd1 vccd1
+ _14059_/X sky130_fd_sc_hd__a221o_1
XFILLER_45_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18936_ _18936_/CLK _18936_/D vssd1 vssd1 vccd1 vccd1 _18936_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_113_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18867_ _18870_/CLK _18867_/D vssd1 vssd1 vccd1 vccd1 _18867_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_39_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17818_ _17821_/CLK _17818_/D vssd1 vssd1 vccd1 vccd1 _17818_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_95_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19062__33 vssd1 vssd1 vccd1 vccd1 _19062__33/HI _19156_/A sky130_fd_sc_hd__conb_1
XFILLER_67_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18798_ _18811_/CLK _18798_/D vssd1 vssd1 vccd1 vccd1 _18798_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_94_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17749_ _17749_/A vssd1 vssd1 vccd1 vccd1 _19017_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_54_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_240 _18358_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_251 _09103_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_262 _14030_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_165_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_273 _18889_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_195_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09103_ _09103_/A _09103_/B _09103_/C _09103_/D vssd1 vssd1 vccd1 vccd1 _09104_/C
+ sky130_fd_sc_hd__and4_1
XFILLER_202_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09034_ _09034_/A vssd1 vssd1 vccd1 vccd1 _09034_/Y sky130_fd_sc_hd__inv_2
XFILLER_190_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_144_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_172_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_104_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09936_ _09418_/A _09413_/D _09408_/D _09418_/C _09959_/A _09935_/X vssd1 vssd1 vccd1
+ vccd1 _09936_/X sky130_fd_sc_hd__mux4_1
XFILLER_217_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_219_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_213_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09867_ _09867_/A _09867_/B vssd1 vssd1 vccd1 vccd1 _09868_/B sky130_fd_sc_hd__nand2_1
XTAP_691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_213_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_93_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09798_ _09813_/A _09795_/Y _09817_/B _09797_/Y vssd1 vssd1 vccd1 vccd1 _09810_/C
+ sky130_fd_sc_hd__a211o_1
XTAP_3237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11760_ _11761_/A _11760_/B vssd1 vssd1 vccd1 vccd1 _11763_/A sky130_fd_sc_hd__nand2_1
XTAP_2558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_148_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10711_ _10790_/B vssd1 vssd1 vccd1 vccd1 _10805_/B sky130_fd_sc_hd__buf_2
XFILLER_13_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11691_ _17852_/Q _11706_/A vssd1 vssd1 vccd1 vccd1 _11691_/Y sky130_fd_sc_hd__nand2_1
XFILLER_41_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_224_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10642_ _10810_/S vssd1 vssd1 vccd1 vccd1 _10737_/S sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_139_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13430_ _11937_/C _13426_/Y _13422_/Y _13429_/Y _11396_/B vssd1 vssd1 vccd1 vccd1
+ _13430_/X sky130_fd_sc_hd__o32a_1
XFILLER_179_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_220_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_224_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13361_ _18105_/Q _13356_/Y _17705_/S vssd1 vssd1 vccd1 vccd1 _13362_/A sky130_fd_sc_hd__mux2_1
XFILLER_210_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10573_ _09314_/B _09319_/A _09319_/C _09309_/C _09688_/A _10036_/X vssd1 vssd1 vccd1
+ vccd1 _10573_/X sky130_fd_sc_hd__mux4_2
XFILLER_127_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_220_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15100_ _18400_/Q _18364_/Q _15100_/S vssd1 vssd1 vccd1 vccd1 _15100_/X sky130_fd_sc_hd__mux2_1
XFILLER_177_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12312_ _12312_/A vssd1 vssd1 vccd1 vccd1 _17878_/D sky130_fd_sc_hd__clkbuf_1
X_16080_ _18632_/Q _18596_/Q _16091_/S vssd1 vssd1 vccd1 vccd1 _16080_/X sky130_fd_sc_hd__mux2_1
XFILLER_154_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13292_ _13292_/A _13292_/B _13292_/C _13292_/D vssd1 vssd1 vccd1 vccd1 _13311_/A
+ sky130_fd_sc_hd__or4_2
XFILLER_166_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_181_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15031_ _15042_/A _15175_/B _15054_/C vssd1 vssd1 vccd1 vccd1 _15031_/X sky130_fd_sc_hd__or3_1
X_12243_ _11648_/X _12242_/X _12269_/B vssd1 vssd1 vccd1 vccd1 _12243_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_174_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12174_ _17846_/Q _12183_/B vssd1 vssd1 vccd1 vccd1 _12174_/X sky130_fd_sc_hd__and2_1
XFILLER_64_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11125_ _11403_/A vssd1 vssd1 vccd1 vccd1 _11467_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_190_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_231_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16982_ _14357_/X _16975_/X _16978_/X _16981_/Y _14618_/X vssd1 vssd1 vccd1 vccd1
+ _18808_/D sky130_fd_sc_hd__o311a_1
XFILLER_95_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18721_ _18722_/CLK _18721_/D vssd1 vssd1 vccd1 vccd1 _18721_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_114_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15933_ _16566_/A vssd1 vssd1 vccd1 vccd1 _16193_/A sky130_fd_sc_hd__clkbuf_2
XTAP_5140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11056_ _17786_/Q vssd1 vssd1 vccd1 vccd1 _11336_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_231_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10007_ _12065_/A _10007_/B vssd1 vssd1 vccd1 vccd1 _10008_/A sky130_fd_sc_hd__and2b_1
X_18652_ _18663_/CLK _18652_/D vssd1 vssd1 vccd1 vccd1 _18652_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_5184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_231_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15864_ _18581_/Q _18545_/Q _15879_/S vssd1 vssd1 vccd1 vccd1 _15864_/X sky130_fd_sc_hd__mux2_1
XTAP_4450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17603_ _17631_/A vssd1 vssd1 vccd1 vccd1 _17603_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_4483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14815_ _14814_/B _14813_/X _14814_/Y _14799_/X vssd1 vssd1 vccd1 vccd1 _18293_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_97_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18583_ _18590_/CLK _18583_/D vssd1 vssd1 vccd1 vccd1 _18583_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_4494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15795_ _15818_/A _15795_/B vssd1 vssd1 vccd1 vccd1 _15795_/Y sky130_fd_sc_hd__nand2_1
XTAP_3760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17534_ _17544_/A _17534_/B vssd1 vssd1 vccd1 vccd1 _17534_/Y sky130_fd_sc_hd__nand2_1
XTAP_3793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14746_ _14928_/A vssd1 vssd1 vccd1 vccd1 _14793_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_18_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11958_ _11984_/C _11280_/Y _11985_/A _11974_/B vssd1 vssd1 vccd1 vccd1 _11958_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_17_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_1306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17465_ _17509_/A _17469_/B vssd1 vssd1 vccd1 vccd1 _17465_/Y sky130_fd_sc_hd__nand2_1
X_10909_ _10678_/X _12094_/A _10904_/X _10906_/X _10908_/X vssd1 vssd1 vccd1 vccd1
+ _10910_/B sky130_fd_sc_hd__o311a_1
XFILLER_199_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14677_ _16945_/A vssd1 vssd1 vccd1 vccd1 _16949_/A sky130_fd_sc_hd__clkbuf_4
X_11889_ _12207_/A _11889_/B vssd1 vssd1 vccd1 vccd1 _17836_/D sky130_fd_sc_hd__nor2_1
X_19204_ _19204_/A _08971_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[4] sky130_fd_sc_hd__ebufn_8
XFILLER_32_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16416_ _18710_/Q _18674_/Q _16421_/S vssd1 vssd1 vccd1 vccd1 _16416_/X sky130_fd_sc_hd__mux2_1
XFILLER_189_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13628_ _18459_/Q _13588_/A _13861_/A _18474_/Q vssd1 vssd1 vccd1 vccd1 _13628_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_177_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17396_ _17395_/B _17394_/X _17395_/Y _17380_/X vssd1 vssd1 vccd1 vccd1 _18911_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_220_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19135_ _19135_/A _09046_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[5] sky130_fd_sc_hd__ebufn_8
X_16347_ _16353_/B _16345_/X _16346_/X _16334_/X vssd1 vssd1 vccd1 vccd1 _18657_/D
+ sky130_fd_sc_hd__o211a_1
X_13559_ _13559_/A vssd1 vssd1 vccd1 vccd1 _13560_/A sky130_fd_sc_hd__buf_4
XFILLER_34_1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16278_ _17222_/A vssd1 vssd1 vccd1 vccd1 _16521_/A sky130_fd_sc_hd__buf_2
XFILLER_172_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18017_ _18224_/CLK _18017_/D vssd1 vssd1 vccd1 vccd1 _18017_/Q sky130_fd_sc_hd__dfxtp_1
X_15229_ _15229_/A _15229_/B vssd1 vssd1 vccd1 vccd1 _15239_/B sky130_fd_sc_hd__nor2_2
XFILLER_160_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_126_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09721_ _09657_/X _09691_/X _09711_/X _09718_/X _09720_/X vssd1 vssd1 vccd1 vccd1
+ _09728_/C sky130_fd_sc_hd__a32o_1
XFILLER_41_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18919_ _18959_/CLK _18919_/D vssd1 vssd1 vccd1 vccd1 _18919_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_101_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_228_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_227_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_210_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09652_ _09653_/A _09653_/B vssd1 vssd1 vccd1 vccd1 _09692_/A sky130_fd_sc_hd__nor2_8
XFILLER_83_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_228_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_215_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09583_ _09600_/A _09583_/B vssd1 vssd1 vccd1 vccd1 _09585_/C sky130_fd_sc_hd__xnor2_1
XFILLER_209_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_230_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_223_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_168_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_211_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_192_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09017_ _09029_/A vssd1 vssd1 vccd1 vccd1 _09022_/A sky130_fd_sc_hd__buf_12
XFILLER_163_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_219_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_104_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_132_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09919_ _09919_/A _09919_/B vssd1 vssd1 vccd1 vccd1 _12122_/A sky130_fd_sc_hd__nand2_4
XFILLER_120_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_218_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12930_ _12930_/A vssd1 vssd1 vccd1 vccd1 _12933_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_58_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_219_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_219_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_207_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12861_ _17951_/Q _12865_/C vssd1 vssd1 vccd1 vccd1 _12864_/A sky130_fd_sc_hd__and2_1
XTAP_2311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14600_ _16862_/A vssd1 vssd1 vccd1 vccd1 _16865_/A sky130_fd_sc_hd__buf_6
XFILLER_61_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11812_ _11905_/A _11812_/B _11812_/C vssd1 vssd1 vccd1 vccd1 _11867_/A sky130_fd_sc_hd__and3b_2
XTAP_2344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15580_ _15583_/B _15577_/X _15579_/Y _15575_/X vssd1 vssd1 vccd1 vccd1 _18475_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_27_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12792_ _17961_/Q vssd1 vssd1 vccd1 vccd1 _12792_/X sky130_fd_sc_hd__clkbuf_2
XTAP_2366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14531_ _14598_/A vssd1 vssd1 vccd1 vccd1 _14584_/B sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_1643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11743_ _11732_/A _11732_/B _11742_/X vssd1 vssd1 vccd1 vccd1 _11826_/C sky130_fd_sc_hd__o21a_1
XTAP_1654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_226_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_202_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_183_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_230_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17250_ _17252_/B _17248_/X _17249_/Y _17241_/X vssd1 vssd1 vccd1 vccd1 _18874_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_1687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14462_ _14463_/A _14463_/B _14461_/X _14340_/X vssd1 vssd1 vccd1 vccd1 _18207_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_105_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11674_ _11672_/A _11673_/A _12253_/A _11669_/B _11669_/A vssd1 vssd1 vccd1 vccd1
+ _11674_/X sky130_fd_sc_hd__a311o_1
XFILLER_224_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16201_ _18659_/Q _18623_/Q _16215_/S vssd1 vssd1 vccd1 vccd1 _16201_/X sky130_fd_sc_hd__mux2_1
XFILLER_122_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13413_ _13409_/X _11218_/X _13412_/X _10990_/X _13016_/X vssd1 vssd1 vccd1 vccd1
+ _18151_/D sky130_fd_sc_hd__a32o_1
XFILLER_186_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17181_ _17197_/A vssd1 vssd1 vccd1 vccd1 _17181_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_70_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10625_ _10629_/A _10625_/B vssd1 vssd1 vccd1 vccd1 _10661_/A sky130_fd_sc_hd__xnor2_4
XFILLER_224_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14393_ _18189_/Q _14404_/A _14386_/B vssd1 vssd1 vccd1 vccd1 _14393_/X sky130_fd_sc_hd__a21o_1
XFILLER_195_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16132_ _16132_/A _16132_/B vssd1 vssd1 vccd1 vccd1 _16132_/Y sky130_fd_sc_hd__nand2_1
XFILLER_155_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_183_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10556_ _09181_/D _09176_/D _09186_/A _09181_/A _10542_/A _10464_/X vssd1 vssd1 vccd1
+ vccd1 _10556_/X sky130_fd_sc_hd__mux4_1
X_13344_ _13344_/A vssd1 vssd1 vccd1 vccd1 _13344_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_154_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16063_ _18592_/Q _16064_/B _16062_/Y _16048_/X vssd1 vssd1 vccd1 vccd1 _18592_/D
+ sky130_fd_sc_hd__o211a_1
X_13275_ _19022_/Q _19021_/Q _19024_/Q _19023_/Q vssd1 vssd1 vccd1 vccd1 _13278_/B
+ sky130_fd_sc_hd__or4_1
X_10487_ _10483_/X _10485_/X _11925_/A vssd1 vssd1 vccd1 vccd1 _10487_/X sky130_fd_sc_hd__mux2_1
XFILLER_154_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15014_ _15156_/A _15136_/C vssd1 vssd1 vccd1 vccd1 _15025_/B sky130_fd_sc_hd__nor2_2
XFILLER_29_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12226_ _12221_/Y _12239_/C _12223_/X _12346_/A vssd1 vssd1 vccd1 vccd1 _17855_/D
+ sky130_fd_sc_hd__a211oi_1
XFILLER_155_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12157_ _12158_/A _12158_/B vssd1 vssd1 vccd1 vccd1 _12157_/Y sky130_fd_sc_hd__nand2_1
XFILLER_9_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_151_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11108_ _17797_/Q vssd1 vssd1 vccd1 vccd1 _11359_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_16965_ _16972_/B _16961_/X _16963_/X _16964_/X vssd1 vssd1 vccd1 vccd1 _18804_/D
+ sky130_fd_sc_hd__o211a_1
X_12088_ _12120_/A _12085_/B _12086_/X _12087_/Y vssd1 vssd1 vccd1 vccd1 _12088_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_110_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_209_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18704_ _18708_/CLK _18704_/D vssd1 vssd1 vccd1 vccd1 _18704_/Q sky130_fd_sc_hd__dfxtp_2
X_15916_ _16673_/A vssd1 vssd1 vccd1 vccd1 _16528_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_37_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11039_ _11039_/A vssd1 vssd1 vccd1 vccd1 _17782_/D sky130_fd_sc_hd__clkbuf_1
X_16896_ _17222_/A vssd1 vssd1 vccd1 vccd1 _17164_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_37_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18635_ _18635_/CLK _18635_/D vssd1 vssd1 vccd1 vccd1 _18635_/Q sky130_fd_sc_hd__dfxtp_2
X_15847_ _15857_/A _15997_/B _15870_/C vssd1 vssd1 vccd1 vccd1 _15847_/X sky130_fd_sc_hd__or3_1
XTAP_4280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18566_ _18571_/CLK _18566_/D vssd1 vssd1 vccd1 vccd1 _18566_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_52_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15778_ _18559_/Q _18523_/Q _15790_/S vssd1 vssd1 vccd1 vccd1 _15778_/X sky130_fd_sc_hd__mux2_1
XTAP_3590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17517_ _17517_/A vssd1 vssd1 vccd1 vccd1 _17517_/X sky130_fd_sc_hd__buf_2
X_14729_ _14753_/A _14729_/B vssd1 vssd1 vccd1 vccd1 _14729_/Y sky130_fd_sc_hd__nand2_1
X_18497_ _18497_/CLK _18497_/D vssd1 vssd1 vccd1 vccd1 _18497_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_205_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_221_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17448_ _17448_/A vssd1 vssd1 vccd1 vccd1 _17493_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_178_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17379_ _17392_/A _17383_/B vssd1 vssd1 vccd1 vccd1 _17379_/Y sky130_fd_sc_hd__nand2_1
XFILLER_119_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_9_wb_clk_i clkbuf_5_4_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17933_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_174_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_203_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_1240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_204_wb_clk_i clkbuf_5_6_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18986_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_138_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_173_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_1216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_6 _09114_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_214_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09704_ _09704_/A _09704_/B vssd1 vssd1 vccd1 vccd1 _10568_/A sky130_fd_sc_hd__or2_1
XFILLER_56_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_229_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_228_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_1340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09635_ _09645_/A _09645_/B _09634_/X vssd1 vssd1 vccd1 vccd1 _09637_/B sky130_fd_sc_hd__a21oi_1
XFILLER_216_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_215_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09566_ _09575_/A _09575_/B vssd1 vssd1 vccd1 vccd1 _09576_/B sky130_fd_sc_hd__xnor2_1
XFILLER_93_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_215_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_231_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_180_1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09497_ _18195_/Q _09497_/B vssd1 vssd1 vccd1 vccd1 _09498_/B sky130_fd_sc_hd__or2_1
XFILLER_196_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_180_1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_221_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10410_ _10542_/A vssd1 vssd1 vccd1 vccd1 _10411_/A sky130_fd_sc_hd__buf_4
XFILLER_139_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11390_ _11390_/A vssd1 vssd1 vccd1 vccd1 _11390_/X sky130_fd_sc_hd__buf_2
XFILLER_109_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10341_ _09921_/X _10339_/X _10340_/X _10605_/B vssd1 vssd1 vccd1 vccd1 _10341_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_180_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_125_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_1176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13060_ _13063_/A _13059_/Y _12776_/X vssd1 vssd1 vccd1 vccd1 _13060_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_124_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10272_ _13410_/A _13410_/B _13410_/C _13410_/D vssd1 vssd1 vccd1 vccd1 _13415_/A
+ sky130_fd_sc_hd__or4_2
XFILLER_3_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12011_ _12011_/A vssd1 vssd1 vccd1 vccd1 _12129_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_191_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16750_ _16755_/B _16747_/X _16749_/X _16740_/X vssd1 vssd1 vccd1 vccd1 _18756_/D
+ sky130_fd_sc_hd__o211a_1
X_13962_ _18661_/Q _13714_/X _13698_/A _18652_/Q _13961_/X vssd1 vssd1 vccd1 vccd1
+ _13962_/X sky130_fd_sc_hd__a221o_2
XFILLER_48_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15701_ _15708_/B _15698_/X _15699_/X _15700_/X vssd1 vssd1 vccd1 vccd1 _18504_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_79_wb_clk_i clkbuf_5_23_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18608_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_46_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12913_ _12913_/A _17968_/Q _12913_/C vssd1 vssd1 vccd1 vccd1 _12913_/X sky130_fd_sc_hd__and3_1
XFILLER_98_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_219_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16681_ _16695_/A _16686_/B vssd1 vssd1 vccd1 vccd1 _16681_/Y sky130_fd_sc_hd__nand2_1
XFILLER_19_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13893_ _18595_/Q _13505_/A _13764_/A _18619_/Q vssd1 vssd1 vccd1 vccd1 _13893_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_111_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18420_ _18423_/CLK _18420_/D vssd1 vssd1 vccd1 vccd1 _18420_/Q sky130_fd_sc_hd__dfxtp_4
X_15632_ _18524_/Q _18488_/Q _15642_/S vssd1 vssd1 vccd1 vccd1 _15632_/X sky130_fd_sc_hd__mux2_1
XTAP_2130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12844_ _12844_/A vssd1 vssd1 vccd1 vccd1 _17946_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_222_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18351_ _18356_/CLK _18351_/D vssd1 vssd1 vccd1 vccd1 _18351_/Q sky130_fd_sc_hd__dfxtp_4
XTAP_2174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15563_ _15613_/A _16007_/B _15574_/C vssd1 vssd1 vccd1 vccd1 _15563_/X sky130_fd_sc_hd__or3_1
XFILLER_15_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12775_ _12775_/A _12951_/B vssd1 vssd1 vccd1 vccd1 _12786_/B sky130_fd_sc_hd__nor2_2
XTAP_2196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17302_ _18923_/Q _18887_/Q _17317_/S vssd1 vssd1 vccd1 vccd1 _17302_/X sky130_fd_sc_hd__mux2_1
XFILLER_199_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14514_ _14512_/Y _14513_/X _11822_/X _14372_/B vssd1 vssd1 vccd1 vccd1 _18228_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_202_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18282_ _18290_/CLK _18282_/D vssd1 vssd1 vccd1 vccd1 _18282_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11726_ _11767_/B _11753_/A _12509_/A vssd1 vssd1 vccd1 vccd1 _11726_/Y sky130_fd_sc_hd__o21ai_1
X_15494_ _18490_/Q _18454_/Q _15494_/S vssd1 vssd1 vccd1 vccd1 _15494_/X sky130_fd_sc_hd__mux2_1
XTAP_1495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17233_ _18906_/Q _18870_/Q _17244_/S vssd1 vssd1 vccd1 vccd1 _17233_/X sky130_fd_sc_hd__mux2_1
X_14445_ _18202_/Q _14445_/B vssd1 vssd1 vccd1 vccd1 _14445_/Y sky130_fd_sc_hd__nor2_1
X_11657_ _11681_/C _11305_/X _11595_/Y _11795_/A vssd1 vssd1 vccd1 vccd1 _11658_/A
+ sky130_fd_sc_hd__o22a_1
XFILLER_200_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17164_ _17164_/A vssd1 vssd1 vccd1 vccd1 _17210_/A sky130_fd_sc_hd__buf_2
XFILLER_70_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10608_ _13000_/B _10619_/B vssd1 vssd1 vccd1 vccd1 _10731_/A sky130_fd_sc_hd__xnor2_4
XFILLER_196_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14376_ _18187_/Q _14375_/B _14373_/X vssd1 vssd1 vccd1 vccd1 _14376_/Y sky130_fd_sc_hd__a21oi_1
X_11588_ _13442_/A _13427_/A _13448_/A vssd1 vssd1 vccd1 vccd1 _11588_/X sky130_fd_sc_hd__or3_1
XFILLER_156_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16115_ _16115_/A _16716_/B _16115_/C vssd1 vssd1 vccd1 vccd1 _16115_/X sky130_fd_sc_hd__or3_1
XFILLER_143_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13327_ _13318_/X _13326_/X _13324_/A vssd1 vssd1 vccd1 vccd1 _13327_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_7_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10539_ _09678_/X _09677_/X _09676_/X _10600_/B _10522_/A _10509_/S vssd1 vssd1 vccd1
+ vccd1 _10539_/X sky130_fd_sc_hd__mux4_1
XFILLER_128_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17095_ _17136_/A _17528_/B _17109_/C vssd1 vssd1 vccd1 vccd1 _17095_/X sky130_fd_sc_hd__or3_1
XFILLER_155_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16046_ _16062_/A _16051_/B vssd1 vssd1 vccd1 vccd1 _16046_/Y sky130_fd_sc_hd__nand2_1
XFILLER_115_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13258_ _13266_/A _18083_/Q vssd1 vssd1 vccd1 vccd1 _13259_/A sky130_fd_sc_hd__and2_1
XFILLER_89_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_142_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12209_ _11706_/A _12200_/X _11704_/A vssd1 vssd1 vccd1 vccd1 _12209_/X sky130_fd_sc_hd__a21o_1
X_13189_ _13197_/A _18052_/Q vssd1 vssd1 vccd1 vccd1 _13190_/A sky130_fd_sc_hd__and2_1
XFILLER_36_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_229_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_215_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17997_ _18151_/CLK _17997_/D vssd1 vssd1 vccd1 vccd1 _17997_/Q sky130_fd_sc_hd__dfxtp_1
X_16948_ _17148_/A vssd1 vssd1 vccd1 vccd1 _17015_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_42_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_1282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16879_ _16879_/A vssd1 vssd1 vccd1 vccd1 _16936_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_168_1334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09420_ _09420_/A _09419_/Y vssd1 vssd1 vccd1 vccd1 _09420_/X sky130_fd_sc_hd__or2b_1
X_18618_ _18623_/CLK _18618_/D vssd1 vssd1 vccd1 vccd1 _18618_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_37_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09351_ _18413_/Q _18412_/Q _18411_/Q vssd1 vssd1 vccd1 vccd1 _10389_/A sky130_fd_sc_hd__or3_4
X_18549_ _18557_/CLK _18549_/D vssd1 vssd1 vccd1 vccd1 _18549_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_212_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09282_ _09282_/A _09282_/B _09282_/C _09282_/D vssd1 vssd1 vccd1 vccd1 _09288_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_221_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_118_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_119_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_173_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08997_ _08997_/A vssd1 vssd1 vccd1 vccd1 _08997_/Y sky130_fd_sc_hd__inv_2
XFILLER_87_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_229_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_1238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_1298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_216_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09618_ _18126_/Q _09618_/B vssd1 vssd1 vccd1 vccd1 _09664_/A sky130_fd_sc_hd__xor2_4
XFILLER_189_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_204_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10890_ _09376_/C _09381_/B _09386_/D _09381_/D _10060_/X _10085_/S vssd1 vssd1 vccd1
+ vccd1 _10890_/X sky130_fd_sc_hd__mux4_1
XFILLER_225_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09549_ _18108_/Q _09549_/B vssd1 vssd1 vccd1 vccd1 _09570_/B sky130_fd_sc_hd__xnor2_1
XFILLER_70_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12560_ _17920_/Q vssd1 vssd1 vccd1 vccd1 _12570_/B sky130_fd_sc_hd__clkinv_2
XFILLER_140_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11511_ _11522_/A _11530_/B vssd1 vssd1 vccd1 vccd1 _11512_/C sky130_fd_sc_hd__nor2_1
XFILLER_197_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_197_wb_clk_i _18176_/CLK vssd1 vssd1 vccd1 vccd1 _18178_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_184_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12491_ _12491_/A vssd1 vssd1 vccd1 vccd1 _17909_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_12_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14230_ _14300_/A vssd1 vssd1 vccd1 vccd1 _17709_/B sky130_fd_sc_hd__clkbuf_2
Xclkbuf_leaf_126_wb_clk_i clkbuf_5_25_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18398_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_137_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11442_ _11442_/A _11442_/B vssd1 vssd1 vccd1 vccd1 _11652_/B sky130_fd_sc_hd__nor2_1
XFILLER_7_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_221_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11373_ _11467_/C _11495_/B _11452_/A vssd1 vssd1 vccd1 vccd1 _11374_/B sky130_fd_sc_hd__o21a_1
X_14161_ _18974_/Q _13621_/A _13568_/X _18968_/Q _14160_/X vssd1 vssd1 vccd1 vccd1
+ _14161_/X sky130_fd_sc_hd__a221o_1
XFILLER_166_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13112_ _13118_/A _18017_/Q vssd1 vssd1 vccd1 vccd1 _13113_/A sky130_fd_sc_hd__and2_1
X_10324_ _09248_/A _09243_/A _09253_/B _10097_/A _10294_/X _09971_/S vssd1 vssd1 vccd1
+ vccd1 _10324_/X sky130_fd_sc_hd__mux4_1
X_14092_ _18416_/Q _14019_/X _14030_/X _18440_/Q _14091_/X vssd1 vssd1 vccd1 vccd1
+ _14092_/X sky130_fd_sc_hd__a221o_1
XFILLER_166_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13043_ _13049_/A _13043_/B vssd1 vssd1 vccd1 vccd1 _13044_/A sky130_fd_sc_hd__and2_1
X_17920_ _18988_/CLK _17920_/D vssd1 vssd1 vccd1 vccd1 _17920_/Q sky130_fd_sc_hd__dfxtp_2
X_10255_ _10253_/A _10188_/B _10186_/X vssd1 vssd1 vccd1 vccd1 _11913_/S sky130_fd_sc_hd__a21oi_1
XFILLER_106_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17851_ _17851_/CLK _17851_/D vssd1 vssd1 vccd1 vccd1 _17851_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_67_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10186_ _18100_/Q _10623_/A vssd1 vssd1 vccd1 vccd1 _10186_/X sky130_fd_sc_hd__and2_1
XFILLER_182_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16802_ _18806_/Q _18770_/Q _16802_/S vssd1 vssd1 vccd1 vccd1 _16802_/X sky130_fd_sc_hd__mux2_1
XFILLER_120_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17782_ _18126_/CLK _17782_/D vssd1 vssd1 vccd1 vccd1 _17782_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_226_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14994_ _18374_/Q _18338_/Q _14994_/S vssd1 vssd1 vccd1 vccd1 _14994_/X sky130_fd_sc_hd__mux2_1
XFILLER_59_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_219_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16733_ _18752_/Q _16732_/B _16732_/Y _16724_/X vssd1 vssd1 vccd1 vccd1 _18752_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_75_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13945_ _18790_/Q _13522_/A _13943_/X _13944_/X vssd1 vssd1 vccd1 vccd1 _13945_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_208_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_223_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_228_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16664_ _16727_/A vssd1 vssd1 vccd1 vccd1 _16794_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_61_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13876_ _18898_/Q _13524_/A _13619_/A _18886_/Q vssd1 vssd1 vccd1 vccd1 _13876_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_201_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15615_ _15630_/A _15618_/B vssd1 vssd1 vccd1 vccd1 _15615_/Y sky130_fd_sc_hd__nand2_1
X_18403_ _18432_/CLK _18403_/D vssd1 vssd1 vccd1 vccd1 _18403_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_90_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12827_ _17939_/Q _17968_/Q vssd1 vssd1 vccd1 vccd1 _12827_/Y sky130_fd_sc_hd__xnor2_1
X_16595_ _18754_/Q _18718_/Q _16598_/S vssd1 vssd1 vccd1 vccd1 _16595_/X sky130_fd_sc_hd__mux2_1
XFILLER_76_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_222_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18334_ _18373_/CLK _18334_/D vssd1 vssd1 vccd1 vccd1 _18334_/Q sky130_fd_sc_hd__dfxtp_2
X_15546_ _15570_/A _15546_/B vssd1 vssd1 vccd1 vccd1 _15546_/Y sky130_fd_sc_hd__nand2_1
XTAP_1270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12758_ _18062_/Q _18036_/Q _12919_/B _12948_/C vssd1 vssd1 vccd1 vccd1 _12758_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_1281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_231_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18265_ _18266_/CLK _18265_/D vssd1 vssd1 vccd1 vccd1 _18265_/Q sky130_fd_sc_hd__dfxtp_1
X_11709_ _17853_/Q _11709_/B _11696_/C vssd1 vssd1 vccd1 vccd1 _11709_/X sky130_fd_sc_hd__or3b_1
XFILLER_37_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15477_ _18145_/Q _15772_/B vssd1 vssd1 vccd1 vccd1 _15589_/A sky130_fd_sc_hd__nand2_4
X_12689_ _12688_/A _12688_/B _12537_/S vssd1 vssd1 vccd1 vccd1 _12689_/X sky130_fd_sc_hd__o21a_1
XFILLER_204_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17216_ _18903_/Q _18867_/Q _17221_/S vssd1 vssd1 vccd1 vccd1 _17216_/X sky130_fd_sc_hd__mux2_1
XFILLER_129_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14428_ _14428_/A vssd1 vssd1 vccd1 vccd1 _14428_/X sky130_fd_sc_hd__clkbuf_2
X_18196_ _18196_/CLK _18196_/D vssd1 vssd1 vccd1 vccd1 _18196_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_200_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17147_ _18885_/Q _18849_/Q _17151_/S vssd1 vssd1 vccd1 vccd1 _17147_/X sky130_fd_sc_hd__mux2_1
XFILLER_143_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14359_ _17943_/Q _14272_/X _14358_/X _12972_/X vssd1 vssd1 vccd1 vccd1 _18183_/D
+ sky130_fd_sc_hd__a211o_1
XFILLER_115_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17078_ _17078_/A vssd1 vssd1 vccd1 vccd1 _17094_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_6_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16029_ _16027_/B _16026_/X _16027_/Y _16028_/X vssd1 vssd1 vccd1 vccd1 _18584_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_170_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_1322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_1366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_226_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_211_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_213_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_214_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09403_ _09403_/A _09403_/B _09403_/C vssd1 vssd1 vccd1 vccd1 _09420_/A sky130_fd_sc_hd__and3_1
XFILLER_25_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09334_ _18527_/Q _18526_/Q _18525_/Q vssd1 vssd1 vccd1 vccd1 _09337_/B sky130_fd_sc_hd__or3_4
XFILLER_55_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_205_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_1367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_179_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09265_ _09265_/A _10813_/A _09265_/C _09265_/D vssd1 vssd1 vccd1 vccd1 _09271_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_21_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09196_ _18572_/Q _18571_/Q _18570_/Q vssd1 vssd1 vccd1 vccd1 _09198_/C sky130_fd_sc_hd__or3_4
XFILLER_154_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_193_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_1260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10040_ _10040_/A vssd1 vssd1 vccd1 vccd1 _10069_/A sky130_fd_sc_hd__clkbuf_4
XTAP_5514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11991_ _12044_/A _13710_/B vssd1 vssd1 vccd1 vccd1 _12102_/B sky130_fd_sc_hd__nand2_2
XFILLER_28_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_217_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13730_ _13730_/A vssd1 vssd1 vccd1 vccd1 _13730_/X sky130_fd_sc_hd__buf_4
XFILLER_216_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10942_ _10942_/A vssd1 vssd1 vccd1 vccd1 _10948_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_16_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_1294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_205_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_1215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13661_ _18957_/Q _13651_/X _13656_/X _13660_/X vssd1 vssd1 vccd1 vccd1 _13661_/X
+ sky130_fd_sc_hd__a211o_1
X_10873_ _10859_/S _10870_/X _10872_/X _10838_/A vssd1 vssd1 vccd1 vccd1 _10873_/X
+ sky130_fd_sc_hd__a211o_1
X_15400_ _15442_/A _15403_/B vssd1 vssd1 vccd1 vccd1 _15400_/Y sky130_fd_sc_hd__nand2_1
XFILLER_71_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12612_ _12612_/A _12612_/B vssd1 vssd1 vccd1 vccd1 _12613_/B sky130_fd_sc_hd__xnor2_1
X_16380_ _16672_/A _16504_/C vssd1 vssd1 vccd1 vccd1 _16392_/B sky130_fd_sc_hd__nor2_2
XPHY_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_213_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13592_ _13592_/A vssd1 vssd1 vccd1 vccd1 _13592_/X sky130_fd_sc_hd__buf_6
XPHY_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15331_ _16839_/A vssd1 vssd1 vccd1 vccd1 _15935_/B sky130_fd_sc_hd__buf_2
XPHY_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12543_ _17920_/Q _17917_/Q vssd1 vssd1 vccd1 vccd1 _12543_/X sky130_fd_sc_hd__and2b_1
XPHY_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_223_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18050_ _18052_/CLK _18050_/D vssd1 vssd1 vccd1 vccd1 _18050_/Q sky130_fd_sc_hd__dfxtp_1
X_15262_ _18440_/Q _18404_/Q _15267_/S vssd1 vssd1 vccd1 vccd1 _15262_/X sky130_fd_sc_hd__mux2_1
XFILLER_12_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12474_ _17907_/Q _12499_/C vssd1 vssd1 vccd1 vccd1 _12475_/A sky130_fd_sc_hd__xor2_1
X_17001_ _17435_/A _17109_/C vssd1 vssd1 vccd1 vccd1 _17010_/B sky130_fd_sc_hd__nor2_2
XFILLER_184_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14213_ _18210_/Q _18209_/Q _18208_/Q _14233_/A vssd1 vssd1 vccd1 vccd1 _14213_/Y
+ sky130_fd_sc_hd__nor4_1
XFILLER_137_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11425_ _11622_/A _11420_/X _11424_/X vssd1 vssd1 vccd1 vccd1 _11425_/Y sky130_fd_sc_hd__a21oi_1
X_15193_ _18422_/Q _18386_/Q _15198_/S vssd1 vssd1 vccd1 vccd1 _15193_/X sky130_fd_sc_hd__mux2_1
XFILLER_32_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_1216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14144_ _18578_/Q _13848_/X _13858_/A _18569_/Q vssd1 vssd1 vccd1 vccd1 _14144_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_153_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11356_ _11404_/A _11541_/B _11453_/B vssd1 vssd1 vccd1 vccd1 _11365_/B sky130_fd_sc_hd__o21a_1
XFILLER_99_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_113_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10307_ _09165_/A _09170_/D _10307_/S vssd1 vssd1 vccd1 vccd1 _10307_/X sky130_fd_sc_hd__mux2_1
XFILLER_4_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14075_ _18722_/Q _13856_/X _13858_/X _18713_/Q _14074_/X vssd1 vssd1 vccd1 vccd1
+ _14075_/X sky130_fd_sc_hd__a221o_1
X_18952_ _18953_/CLK _18952_/D vssd1 vssd1 vccd1 vccd1 _18952_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_3_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11287_ _11287_/A vssd1 vssd1 vccd1 vccd1 _11541_/B sky130_fd_sc_hd__clkbuf_2
Xclkbuf_leaf_94_wb_clk_i _18254_/CLK vssd1 vssd1 vccd1 vccd1 _18266_/CLK sky130_fd_sc_hd__clkbuf_16
X_17903_ _17907_/CLK _17903_/D vssd1 vssd1 vccd1 vccd1 _17903_/Q sky130_fd_sc_hd__dfxtp_1
X_13026_ _17986_/Q _13036_/B vssd1 vssd1 vccd1 vccd1 _13026_/X sky130_fd_sc_hd__or2_1
XFILLER_79_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10238_ _10238_/A _10238_/B vssd1 vssd1 vccd1 vccd1 _10466_/A sky130_fd_sc_hd__xor2_1
XFILLER_117_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18883_ _18907_/CLK _18883_/D vssd1 vssd1 vccd1 vccd1 _18883_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_39_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_230_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_23_wb_clk_i clkbuf_5_4_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18203_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_17834_ _18209_/CLK _17834_/D vssd1 vssd1 vccd1 vccd1 _17834_/Q sky130_fd_sc_hd__dfxtp_1
X_10169_ _10169_/A _10169_/B vssd1 vssd1 vccd1 vccd1 _10170_/B sky130_fd_sc_hd__xor2_1
XFILLER_66_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_208_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14977_ _14977_/A vssd1 vssd1 vccd1 vccd1 _14994_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_130_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17765_ _17765_/A vssd1 vssd1 vccd1 vccd1 _19025_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_66_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_212_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16716_ _16736_/A _16716_/B _16716_/C vssd1 vssd1 vccd1 vccd1 _16716_/X sky130_fd_sc_hd__or3_1
X_13928_ _18250_/Q _13594_/A _13725_/X _18232_/Q vssd1 vssd1 vccd1 vccd1 _13928_/X
+ sky130_fd_sc_hd__a22o_1
X_17696_ _17712_/A _17696_/B vssd1 vssd1 vccd1 vccd1 _17697_/A sky130_fd_sc_hd__and2_1
XFILLER_223_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16647_ _16832_/A vssd1 vssd1 vccd1 vccd1 _16699_/A sky130_fd_sc_hd__clkbuf_2
X_13859_ _18823_/Q _13702_/A _13842_/A _18817_/Q vssd1 vssd1 vccd1 vccd1 _13859_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_23_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_222_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16578_ _16578_/A vssd1 vssd1 vccd1 vccd1 _16628_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_210_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_222_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15529_ _15529_/A vssd1 vssd1 vccd1 vccd1 _15574_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_18317_ _18317_/CLK _18317_/D vssd1 vssd1 vccd1 vccd1 _18317_/Q sky130_fd_sc_hd__dfxtp_4
X_09050_ _09052_/A vssd1 vssd1 vccd1 vccd1 _09050_/Y sky130_fd_sc_hd__inv_2
XFILLER_198_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18248_ _18809_/CLK _18248_/D vssd1 vssd1 vccd1 vccd1 _18248_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_176_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_1310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_1204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_190_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18179_ _18184_/CLK _18179_/D vssd1 vssd1 vccd1 vccd1 _18179_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09952_ _09952_/A _10391_/B vssd1 vssd1 vccd1 vccd1 _09952_/X sky130_fd_sc_hd__or2_1
XFILLER_98_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_106_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09883_ _09882_/A _09883_/B vssd1 vssd1 vccd1 vccd1 _09883_/X sky130_fd_sc_hd__and2b_1
XTAP_851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_85_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_213_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_214_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_207_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_198_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_202_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09317_ _18482_/Q _18481_/Q _18480_/Q vssd1 vssd1 vccd1 vccd1 _09319_/C sky130_fd_sc_hd__or3_2
XFILLER_142_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_220_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_210_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09248_ _09248_/A _09248_/B _09248_/C _10097_/A vssd1 vssd1 vccd1 vccd1 _09254_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_107_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_154_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09179_ _18608_/Q _18607_/Q _18606_/Q vssd1 vssd1 vccd1 vccd1 _09181_/C sky130_fd_sc_hd__or3_4
XFILLER_166_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_108_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11210_ _11210_/A _11210_/B _11210_/C vssd1 vssd1 vccd1 vccd1 _11211_/A sky130_fd_sc_hd__and3_1
XFILLER_108_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12190_ _12499_/C vssd1 vssd1 vccd1 vccd1 _12493_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_218_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_190_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11141_ _13485_/A vssd1 vssd1 vccd1 vccd1 _11795_/A sky130_fd_sc_hd__buf_2
XTAP_6001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_6034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11072_ _11070_/X _17818_/Q _11091_/S vssd1 vssd1 vccd1 vccd1 _11073_/A sky130_fd_sc_hd__mux2_1
XTAP_6045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_1290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14900_ _14935_/A _14900_/B vssd1 vssd1 vccd1 vccd1 _14900_/Y sky130_fd_sc_hd__nand2_1
X_10023_ _10103_/B vssd1 vssd1 vccd1 vccd1 _10956_/B sky130_fd_sc_hd__buf_4
XFILLER_0_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15880_ _15921_/A _16032_/B _15894_/C vssd1 vssd1 vccd1 vccd1 _15880_/X sky130_fd_sc_hd__or3_1
XTAP_4610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14831_ _14856_/A _15268_/B _14843_/C vssd1 vssd1 vccd1 vccd1 _14831_/X sky130_fd_sc_hd__or3_1
XTAP_4654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17550_ _17581_/A vssd1 vssd1 vccd1 vccd1 _17675_/A sky130_fd_sc_hd__clkbuf_1
XTAP_4698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14762_ _14944_/A vssd1 vssd1 vccd1 vccd1 _14810_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_17_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11974_ _12041_/A _11974_/B vssd1 vssd1 vccd1 vccd1 _11980_/A sky130_fd_sc_hd__nor2_1
XTAP_3975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16501_ _16794_/A _16501_/B vssd1 vssd1 vccd1 vccd1 _16510_/B sky130_fd_sc_hd__nor2_1
XFILLER_186_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13713_ _13758_/A vssd1 vssd1 vccd1 vccd1 _13730_/A sky130_fd_sc_hd__clkbuf_4
XTAP_3986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10925_ _09332_/C _09337_/D _09337_/A _09327_/D _10509_/S _10522_/X vssd1 vssd1 vccd1
+ vccd1 _10926_/B sky130_fd_sc_hd__mux4_2
XTAP_3997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17481_ _17519_/A vssd1 vssd1 vccd1 vccd1 _17495_/S sky130_fd_sc_hd__clkbuf_2
X_14693_ _18264_/Q _14700_/B _14690_/X _14692_/X vssd1 vssd1 vccd1 vccd1 _18264_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_16_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_204_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_189_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16432_ _17037_/A _16504_/C vssd1 vssd1 vccd1 vccd1 _16439_/B sky130_fd_sc_hd__nor2_2
X_19220_ _19220_/A _08960_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[20] sky130_fd_sc_hd__ebufn_8
XFILLER_108_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_141_wb_clk_i clkbuf_5_26_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18312_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_13644_ _18897_/Q _13596_/A _13630_/A _18879_/Q vssd1 vssd1 vccd1 vccd1 _13644_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_72_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10856_ _10854_/X _10855_/X _10856_/S vssd1 vssd1 vccd1 vccd1 _10856_/X sky130_fd_sc_hd__mux2_1
XFILLER_31_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_213_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19151_ _19151_/A _09033_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[21] sky130_fd_sc_hd__ebufn_8
XFILLER_198_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16363_ _18698_/Q _18662_/Q _16363_/S vssd1 vssd1 vccd1 vccd1 _16363_/X sky130_fd_sc_hd__mux2_1
XFILLER_125_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_160_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13575_ _13575_/A vssd1 vssd1 vccd1 vccd1 _13575_/X sky130_fd_sc_hd__buf_2
XFILLER_31_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10787_ _10779_/X _10780_/X _10784_/X _10910_/D vssd1 vssd1 vccd1 vccd1 _10787_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_158_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18102_ _18102_/CLK _18102_/D vssd1 vssd1 vccd1 vccd1 _18102_/Q sky130_fd_sc_hd__dfxtp_2
XPHY_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15314_ _15739_/A vssd1 vssd1 vccd1 vccd1 _15404_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_13_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12526_ _13357_/B vssd1 vssd1 vccd1 vccd1 _16673_/A sky130_fd_sc_hd__buf_4
X_16294_ _16329_/A _16294_/B vssd1 vssd1 vccd1 vccd1 _16294_/Y sky130_fd_sc_hd__nand2_1
XFILLER_185_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_184_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18033_ _18035_/CLK _18033_/D vssd1 vssd1 vccd1 vccd1 _18033_/Q sky130_fd_sc_hd__dfxtp_1
X_15245_ _15253_/B _15242_/X _15243_/X _15244_/X vssd1 vssd1 vccd1 vccd1 _18399_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_172_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12457_ _12458_/A _12477_/A _12477_/B vssd1 vssd1 vccd1 vccd1 _12459_/B sky130_fd_sc_hd__a21o_1
X_11408_ _11498_/A _11453_/A vssd1 vssd1 vccd1 vccd1 _11609_/A sky130_fd_sc_hd__nand2_2
X_15176_ _15182_/B _15173_/X _15175_/X _15166_/X vssd1 vssd1 vccd1 vccd1 _18381_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_172_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12388_ _12388_/A _12388_/B _12388_/C vssd1 vssd1 vccd1 vccd1 _12389_/C sky130_fd_sc_hd__or3_1
XFILLER_153_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14127_ _18887_/Q _14017_/X _14122_/X _14126_/X vssd1 vssd1 vccd1 vccd1 _14127_/X
+ sky130_fd_sc_hd__a211o_1
X_11339_ _17877_/Q _11339_/B _11339_/C _11339_/D vssd1 vssd1 vccd1 vccd1 _11339_/Y
+ sky130_fd_sc_hd__nand4_1
XFILLER_207_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14058_ _18392_/Q _13877_/A _13582_/A _18386_/Q vssd1 vssd1 vccd1 vccd1 _14058_/X
+ sky130_fd_sc_hd__a22o_1
X_18935_ _18936_/CLK _18935_/D vssd1 vssd1 vccd1 vccd1 _18935_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_80_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13009_ _13009_/A _13009_/B vssd1 vssd1 vccd1 vccd1 _13009_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_79_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18866_ _18866_/CLK _18866_/D vssd1 vssd1 vccd1 vccd1 _18866_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_39_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_227_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17817_ _17817_/CLK _17817_/D vssd1 vssd1 vccd1 vccd1 _17817_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_82_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18797_ _18811_/CLK _18797_/D vssd1 vssd1 vccd1 vccd1 _18797_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_55_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_229_wb_clk_i _17864_/CLK vssd1 vssd1 vccd1 vccd1 _19034_/CLK sky130_fd_sc_hd__clkbuf_16
X_17748_ _17756_/A _19018_/Q vssd1 vssd1 vccd1 vccd1 _17749_/A sky130_fd_sc_hd__and2_1
XFILLER_130_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_230 _15243_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17679_ _17679_/A vssd1 vssd1 vccd1 vccd1 _18981_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_165_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_241 _18368_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_252 _09109_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_263 _17575_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_211_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XINSDIODE2_274 _18182_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09102_ _18779_/Q _18778_/Q _18777_/Q vssd1 vssd1 vccd1 vccd1 _09103_/D sky130_fd_sc_hd__or3_4
XFILLER_206_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09033_ _09034_/A vssd1 vssd1 vccd1 vccd1 _09033_/Y sky130_fd_sc_hd__inv_2
XFILLER_164_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_176_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_176_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09935_ _10316_/S vssd1 vssd1 vccd1 vccd1 _09935_/X sky130_fd_sc_hd__buf_6
XFILLER_131_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_219_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09866_ _09866_/A _09866_/B vssd1 vssd1 vccd1 vccd1 _09874_/A sky130_fd_sc_hd__xor2_4
XFILLER_218_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_213_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09797_ _09812_/A _09812_/B vssd1 vssd1 vccd1 vccd1 _09797_/Y sky130_fd_sc_hd__nor2_1
XTAP_3216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_1280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10710_ _10731_/A _10710_/B vssd1 vssd1 vccd1 vccd1 _10790_/B sky130_fd_sc_hd__nor2_2
XTAP_1858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11690_ _17851_/Q _17850_/Q vssd1 vssd1 vccd1 vccd1 _11706_/A sky130_fd_sc_hd__and2_1
XFILLER_13_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_201_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10641_ _10716_/A vssd1 vssd1 vccd1 vccd1 _10810_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_224_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_220_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13360_ _14384_/B _13363_/B vssd1 vssd1 vccd1 vccd1 _17705_/S sky130_fd_sc_hd__and2_2
XFILLER_224_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_220_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10572_ _10076_/S _10566_/X _10571_/X _10069_/A vssd1 vssd1 vccd1 vccd1 _10572_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_10_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_167_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12311_ _14504_/B _12333_/C _12311_/C vssd1 vssd1 vccd1 vccd1 _12312_/A sky130_fd_sc_hd__and3_1
X_19108__79 vssd1 vssd1 vccd1 vccd1 _19108__79/HI _19216_/A sky130_fd_sc_hd__conb_1
XFILLER_181_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13291_ _13291_/A _13291_/B _13291_/C _13291_/D vssd1 vssd1 vccd1 vccd1 _13292_/D
+ sky130_fd_sc_hd__or4_1
XFILLER_33_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_182_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15030_ _18381_/Q _18345_/Q _15033_/S vssd1 vssd1 vccd1 vccd1 _15030_/X sky130_fd_sc_hd__mux2_1
X_12242_ _17863_/Q _11642_/X _17864_/Q vssd1 vssd1 vccd1 vccd1 _12242_/X sky130_fd_sc_hd__a21o_1
XFILLER_194_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12173_ _12171_/X _12172_/X _12163_/X vssd1 vssd1 vccd1 vccd1 _17845_/D sky130_fd_sc_hd__o21a_1
XFILLER_218_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_1358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11124_ _17799_/Q vssd1 vssd1 vccd1 vccd1 _11403_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_1_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16981_ _16975_/A _16978_/X _18808_/Q vssd1 vssd1 vccd1 vccd1 _16981_/Y sky130_fd_sc_hd__o21bai_1
XFILLER_77_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18720_ _18722_/CLK _18720_/D vssd1 vssd1 vccd1 vccd1 _18720_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_150_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15932_ _18597_/Q _18561_/Q _15937_/S vssd1 vssd1 vccd1 vccd1 _15932_/X sky130_fd_sc_hd__mux2_1
XTAP_5130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11055_ _11055_/A vssd1 vssd1 vccd1 vccd1 _17785_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_110_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_231_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10006_ _09683_/X _10003_/X _10005_/X _10962_/A vssd1 vssd1 vccd1 vccd1 _10006_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_37_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18651_ _18663_/CLK _18651_/D vssd1 vssd1 vccd1 vccd1 _18651_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_5174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15863_ _15863_/A vssd1 vssd1 vccd1 vccd1 _15879_/S sky130_fd_sc_hd__clkbuf_2
XTAP_5185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14814_ _14814_/A _14814_/B vssd1 vssd1 vccd1 vccd1 _14814_/Y sky130_fd_sc_hd__nand2_1
X_17602_ _17602_/A _17663_/A vssd1 vssd1 vccd1 vccd1 _17602_/Y sky130_fd_sc_hd__nor2_2
XFILLER_97_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_224_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15794_ _18563_/Q _18527_/Q _15809_/S vssd1 vssd1 vccd1 vccd1 _15794_/X sky130_fd_sc_hd__mux2_1
X_18582_ _18582_/CLK _18582_/D vssd1 vssd1 vccd1 vccd1 _18582_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_4484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_205_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14745_ _18312_/Q _18276_/Q _14756_/S vssd1 vssd1 vccd1 vccd1 _14745_/X sky130_fd_sc_hd__mux2_1
XFILLER_51_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17533_ _18983_/Q _18947_/Q _17533_/S vssd1 vssd1 vccd1 vccd1 _17533_/X sky130_fd_sc_hd__mux2_1
XTAP_3794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11957_ _12028_/D _11957_/B vssd1 vssd1 vccd1 vccd1 _11967_/A sky130_fd_sc_hd__or2_1
XFILLER_72_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17464_ _17464_/A vssd1 vssd1 vccd1 vccd1 _17509_/A sky130_fd_sc_hd__buf_2
X_10908_ _10678_/X _10907_/X _10679_/X vssd1 vssd1 vccd1 vccd1 _10908_/X sky130_fd_sc_hd__a21o_1
X_14676_ _14928_/A vssd1 vssd1 vccd1 vccd1 _14734_/A sky130_fd_sc_hd__buf_4
XFILLER_220_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11888_ _18161_/Q _11852_/X _11875_/Y vssd1 vssd1 vccd1 vccd1 _11889_/B sky130_fd_sc_hd__a21oi_1
X_16415_ _16417_/B _16413_/X _16414_/Y _16398_/X vssd1 vssd1 vccd1 vccd1 _18673_/D
+ sky130_fd_sc_hd__o211a_1
X_19203_ _19203_/A _08988_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[3] sky130_fd_sc_hd__ebufn_8
X_13627_ _13703_/A vssd1 vssd1 vccd1 vccd1 _13861_/A sky130_fd_sc_hd__buf_6
X_17395_ _17395_/A _17395_/B vssd1 vssd1 vccd1 vccd1 _17395_/Y sky130_fd_sc_hd__nand2_1
X_10839_ _10867_/A _10834_/X _10836_/X _10838_/X vssd1 vssd1 vccd1 vccd1 _10839_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_158_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16346_ _16371_/A _16785_/B _16358_/C vssd1 vssd1 vccd1 vccd1 _16346_/X sky130_fd_sc_hd__or3_1
XFILLER_186_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19134_ _19134_/A _09049_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[4] sky130_fd_sc_hd__ebufn_8
XFILLER_34_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13558_ _13583_/A vssd1 vssd1 vccd1 vccd1 _13559_/A sky130_fd_sc_hd__buf_6
XFILLER_9_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12509_ _12509_/A _12514_/A vssd1 vssd1 vccd1 vccd1 _12509_/Y sky130_fd_sc_hd__nor2_1
X_16277_ _18676_/Q _18640_/Q _16304_/S vssd1 vssd1 vccd1 vccd1 _16277_/X sky130_fd_sc_hd__mux2_1
X_13489_ _13489_/A vssd1 vssd1 vccd1 vccd1 _13490_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_66_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15228_ _15227_/B _15226_/X _15227_/Y _15224_/X vssd1 vssd1 vccd1 vccd1 _18395_/D
+ sky130_fd_sc_hd__o211a_1
X_18016_ _18224_/CLK _18016_/D vssd1 vssd1 vccd1 vccd1 _18016_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_126_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15159_ _15270_/A vssd1 vssd1 vccd1 vccd1 _15250_/A sky130_fd_sc_hd__buf_2
X_19122__93 vssd1 vssd1 vccd1 vccd1 _19122__93/HI _19230_/A sky130_fd_sc_hd__conb_1
XFILLER_4_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09720_ _09720_/A vssd1 vssd1 vccd1 vccd1 _09720_/X sky130_fd_sc_hd__buf_4
X_18918_ _18927_/CLK _18918_/D vssd1 vssd1 vccd1 vccd1 _18918_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_86_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09651_ _12078_/A _09649_/X _09679_/A vssd1 vssd1 vccd1 vccd1 _09653_/B sky130_fd_sc_hd__a21oi_4
XFILLER_228_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18849_ _18849_/CLK _18849_/D vssd1 vssd1 vccd1 vccd1 _18849_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_95_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_227_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09582_ _09600_/B _09600_/C vssd1 vssd1 vccd1 vccd1 _09583_/B sky130_fd_sc_hd__xor2_1
XFILLER_55_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_215_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_3_7_0_wb_clk_i clkbuf_3_7_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_7_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_223_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_195_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_191_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09016_ _09016_/A vssd1 vssd1 vccd1 vccd1 _09016_/Y sky130_fd_sc_hd__inv_2
XFILLER_3_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_219_1366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09918_ _09918_/A _09918_/B vssd1 vssd1 vccd1 vccd1 _09919_/B sky130_fd_sc_hd__nand2_1
XFILLER_219_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_219_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09849_ _19028_/Q _17973_/Q vssd1 vssd1 vccd1 vccd1 _10627_/B sky130_fd_sc_hd__xor2_4
XFILLER_100_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12860_ _12860_/A vssd1 vssd1 vccd1 vccd1 _17950_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_206_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_227_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11811_ _12041_/A _11282_/B _11832_/B _11281_/A vssd1 vssd1 vccd1 vccd1 _11812_/C
+ sky130_fd_sc_hd__o31ai_1
XTAP_2334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12791_ _17945_/Q vssd1 vssd1 vccd1 vccd1 _12839_/A sky130_fd_sc_hd__inv_2
XTAP_2345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14530_ _17412_/A vssd1 vssd1 vccd1 vccd1 _15150_/B sky130_fd_sc_hd__buf_6
XTAP_1633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11742_ _11742_/A _11742_/B _11742_/C vssd1 vssd1 vccd1 vccd1 _11742_/X sky130_fd_sc_hd__or3_1
XTAP_1644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14461_ _14279_/A _17709_/B _14233_/A vssd1 vssd1 vccd1 vccd1 _14461_/X sky130_fd_sc_hd__a21o_1
XFILLER_109_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11673_ _11673_/A _11673_/B vssd1 vssd1 vccd1 vccd1 _11673_/X sky130_fd_sc_hd__and2_1
XFILLER_41_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16200_ _16202_/B _16198_/X _16199_/Y _16185_/X vssd1 vssd1 vccd1 vccd1 _18622_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_30_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13412_ _13412_/A _13412_/B _13412_/C vssd1 vssd1 vccd1 vccd1 _13412_/X sky130_fd_sc_hd__and3_1
XFILLER_224_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10624_ _18130_/Q _10627_/B _09850_/X vssd1 vssd1 vccd1 vccd1 _10625_/B sky130_fd_sc_hd__a21oi_2
X_17180_ _17213_/A _17180_/B vssd1 vssd1 vccd1 vccd1 _17180_/Y sky130_fd_sc_hd__nand2_1
XFILLER_122_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14392_ _14422_/A vssd1 vssd1 vccd1 vccd1 _14404_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_183_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16131_ _18607_/Q _16132_/B _16130_/Y _16120_/X vssd1 vssd1 vccd1 vccd1 _18607_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_31_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_122_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13343_ _18098_/Q _13336_/X _13342_/X _13339_/X vssd1 vssd1 vccd1 vccd1 _18098_/D
+ sky130_fd_sc_hd__o211a_1
X_10555_ _10555_/A _10555_/B vssd1 vssd1 vccd1 vccd1 _10555_/X sky130_fd_sc_hd__or2_1
XFILLER_183_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16062_ _16062_/A _16064_/B vssd1 vssd1 vccd1 vccd1 _16062_/Y sky130_fd_sc_hd__nand2_1
XFILLER_143_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13274_ _19014_/Q _19013_/Q _19016_/Q _19015_/Q vssd1 vssd1 vccd1 vccd1 _13278_/A
+ sky130_fd_sc_hd__or4_1
XFILLER_108_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10486_ _10926_/A vssd1 vssd1 vccd1 vccd1 _11925_/A sky130_fd_sc_hd__buf_2
X_15013_ _18341_/Q _15012_/B _15012_/Y _15004_/X vssd1 vssd1 vccd1 vccd1 _18341_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_155_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12225_ _12708_/A vssd1 vssd1 vccd1 vccd1 _12346_/A sky130_fd_sc_hd__buf_8
XFILLER_135_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12156_ _12169_/A _12169_/B vssd1 vssd1 vccd1 vccd1 _12158_/B sky130_fd_sc_hd__xnor2_1
XFILLER_155_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_1330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11107_ _11107_/A vssd1 vssd1 vccd1 vccd1 _17796_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_110_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_231_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16964_ _16999_/A vssd1 vssd1 vccd1 vccd1 _16964_/X sky130_fd_sc_hd__clkbuf_2
X_12087_ _14317_/B _12133_/B vssd1 vssd1 vccd1 vccd1 _12087_/Y sky130_fd_sc_hd__nand2_1
XFILLER_1_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18703_ _18708_/CLK _18703_/D vssd1 vssd1 vccd1 vccd1 _18703_/Q sky130_fd_sc_hd__dfxtp_2
X_15915_ _15915_/A _16043_/C vssd1 vssd1 vccd1 vccd1 _15928_/B sky130_fd_sc_hd__nor2_1
X_11038_ _11038_/A _13398_/A _13367_/A _13370_/B vssd1 vssd1 vccd1 vccd1 _11039_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_231_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16895_ _18826_/Q _18790_/Q _16900_/S vssd1 vssd1 vccd1 vccd1 _16895_/X sky130_fd_sc_hd__mux2_1
XFILLER_42_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18634_ _18635_/CLK _18634_/D vssd1 vssd1 vccd1 vccd1 _18634_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_209_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15846_ _18576_/Q _18540_/Q _15859_/S vssd1 vssd1 vccd1 vccd1 _15846_/X sky130_fd_sc_hd__mux2_1
XTAP_4270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_225_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18565_ _18607_/CLK _18565_/D vssd1 vssd1 vccd1 vccd1 _18565_/Q sky130_fd_sc_hd__dfxtp_4
X_15777_ _15782_/B _15775_/X _15776_/X _15763_/X vssd1 vssd1 vccd1 vccd1 _18522_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_3580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12989_ _12989_/A vssd1 vssd1 vccd1 vccd1 _13007_/B sky130_fd_sc_hd__clkbuf_2
XTAP_3591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17516_ _17538_/A _17516_/B _17516_/C vssd1 vssd1 vccd1 vccd1 _17516_/X sky130_fd_sc_hd__or3_1
X_14728_ _18308_/Q _18272_/Q _14736_/S vssd1 vssd1 vccd1 vccd1 _14728_/X sky130_fd_sc_hd__mux2_1
X_18496_ _18496_/CLK _18496_/D vssd1 vssd1 vccd1 vccd1 _18496_/Q sky130_fd_sc_hd__dfxtp_4
XTAP_2890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_220_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14659_ _18257_/Q _14658_/B _14658_/Y _14647_/X vssd1 vssd1 vccd1 vccd1 _18257_/D
+ sky130_fd_sc_hd__o211a_1
X_17447_ _18960_/Q _18924_/Q _17447_/S vssd1 vssd1 vccd1 vccd1 _17447_/X sky130_fd_sc_hd__mux2_1
XFILLER_60_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_220_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_207_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17378_ _18943_/Q _18907_/Q _17386_/S vssd1 vssd1 vccd1 vccd1 _17378_/X sky130_fd_sc_hd__mux2_1
XFILLER_192_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_146_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16329_ _16329_/A _16329_/B vssd1 vssd1 vccd1 vccd1 _16329_/Y sky130_fd_sc_hd__nand2_1
XFILLER_145_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_1277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_7 _10728_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_214_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_228_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09703_ _09703_/A vssd1 vssd1 vccd1 vccd1 _10942_/A sky130_fd_sc_hd__buf_4
XFILLER_56_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_214_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09634_ _18098_/Q _12946_/A vssd1 vssd1 vccd1 vccd1 _09634_/X sky130_fd_sc_hd__and2_1
XFILLER_167_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_215_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09565_ _09565_/A _09565_/B vssd1 vssd1 vccd1 vccd1 _09575_/B sky130_fd_sc_hd__xnor2_1
XFILLER_110_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_212_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_230_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09496_ _18194_/Q _18193_/Q _14409_/B vssd1 vssd1 vccd1 vccd1 _09497_/B sky130_fd_sc_hd__or3_1
XFILLER_93_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_223_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_1368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_221_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_221_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_221_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10340_ _09126_/C _09131_/B _09136_/D _09131_/D _09909_/X _12121_/A vssd1 vssd1 vccd1
+ vccd1 _10340_/X sky130_fd_sc_hd__mux4_1
XFILLER_191_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_191_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_178_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10271_ _10939_/A _10271_/B _10271_/C vssd1 vssd1 vccd1 vccd1 _13410_/D sky130_fd_sc_hd__and3_1
XFILLER_155_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12010_ _12019_/A _11967_/A _12043_/A _12010_/D vssd1 vssd1 vccd1 vccd1 _12011_/A
+ sky130_fd_sc_hd__and4bb_1
XFILLER_151_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_219_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13961_ _18634_/Q _13749_/X _13957_/X _13960_/X vssd1 vssd1 vccd1 vccd1 _13961_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_59_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15700_ _15720_/A vssd1 vssd1 vccd1 vccd1 _15700_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_24_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12912_ _12913_/A _12913_/C _12911_/Y vssd1 vssd1 vccd1 vccd1 _17967_/D sky130_fd_sc_hd__a21oi_1
X_16680_ _18775_/Q _18739_/Q _16694_/S vssd1 vssd1 vccd1 vccd1 _16680_/X sky130_fd_sc_hd__mux2_1
XFILLER_150_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_1262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13892_ _18607_/Q _13666_/X _13624_/A _18601_/Q _13891_/X vssd1 vssd1 vccd1 vccd1
+ _13892_/X sky130_fd_sc_hd__a221o_1
XFILLER_0_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15631_ _15633_/B _15629_/X _15630_/Y _15616_/X vssd1 vssd1 vccd1 vccd1 _18487_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_185_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12843_ _12888_/B _12843_/B _12846_/B vssd1 vssd1 vccd1 vccd1 _12844_/A sky130_fd_sc_hd__and3_1
XTAP_2131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15562_ _15562_/A vssd1 vssd1 vccd1 vccd1 _15613_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_18350_ _18350_/CLK _18350_/D vssd1 vssd1 vccd1 vccd1 _18350_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_61_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12774_ _18152_/Q _12781_/B vssd1 vssd1 vccd1 vccd1 _12951_/B sky130_fd_sc_hd__or2_1
XTAP_2175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14513_ _14515_/B _14513_/B vssd1 vssd1 vccd1 vccd1 _14513_/X sky130_fd_sc_hd__and2_1
X_17301_ _17370_/A vssd1 vssd1 vccd1 vccd1 _17317_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_159_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_48_wb_clk_i clkbuf_5_5_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18858_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_1474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11725_ _11737_/B vssd1 vssd1 vccd1 vccd1 _12509_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_15493_ _15500_/B _15491_/X _15492_/X _15474_/X vssd1 vssd1 vccd1 vccd1 _18453_/D
+ sky130_fd_sc_hd__o211a_1
X_18281_ _18290_/CLK _18281_/D vssd1 vssd1 vccd1 vccd1 _18281_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_14_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_202_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14444_ _14452_/A _14444_/B vssd1 vssd1 vccd1 vccd1 _18201_/D sky130_fd_sc_hd__nor2_1
X_17232_ _17514_/A _17254_/B vssd1 vssd1 vccd1 vccd1 _17240_/B sky130_fd_sc_hd__nor2_2
XFILLER_175_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11656_ _11748_/C _11656_/B vssd1 vssd1 vccd1 vccd1 _11669_/A sky130_fd_sc_hd__nand2_1
XFILLER_128_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10607_ _18129_/Q _10611_/B _09757_/X vssd1 vssd1 vccd1 vccd1 _10619_/B sky130_fd_sc_hd__a21oi_4
X_17163_ _18889_/Q _18853_/Q _17172_/S vssd1 vssd1 vccd1 vccd1 _17163_/X sky130_fd_sc_hd__mux2_1
XFILLER_127_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14375_ _18187_/Q _14375_/B vssd1 vssd1 vccd1 vccd1 _14375_/X sky130_fd_sc_hd__or2_1
XFILLER_128_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11587_ _11780_/A _11783_/A _11587_/C _11586_/X vssd1 vssd1 vccd1 vccd1 _11808_/B
+ sky130_fd_sc_hd__or4b_4
XFILLER_200_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16114_ _16865_/A vssd1 vssd1 vccd1 vccd1 _16716_/B sky130_fd_sc_hd__buf_4
XFILLER_122_1176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13326_ _18093_/Q _13329_/B vssd1 vssd1 vccd1 vccd1 _13326_/X sky130_fd_sc_hd__xor2_1
X_17094_ _18873_/Q _18837_/Q _17094_/S vssd1 vssd1 vccd1 vccd1 _17094_/X sky130_fd_sc_hd__mux2_1
XFILLER_6_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10538_ _10555_/A _10538_/B vssd1 vssd1 vccd1 vccd1 _10538_/X sky130_fd_sc_hd__and2_1
XFILLER_127_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16045_ _18625_/Q _18589_/Q _16050_/S vssd1 vssd1 vccd1 vccd1 _16045_/X sky130_fd_sc_hd__mux2_1
X_13257_ _13257_/A vssd1 vssd1 vccd1 vccd1 _13266_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_142_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10469_ _09237_/A _09227_/B _09232_/C _09237_/C _10464_/X _10235_/A vssd1 vssd1 vccd1
+ vccd1 _10469_/X sky130_fd_sc_hd__mux4_1
XFILLER_89_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12208_ _12444_/B _12358_/B vssd1 vssd1 vccd1 vccd1 _12210_/A sky130_fd_sc_hd__or2_1
XFILLER_130_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13188_ _13199_/A vssd1 vssd1 vccd1 vccd1 _13197_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_96_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12139_ _12139_/A vssd1 vssd1 vccd1 vccd1 _12169_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_111_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17996_ _18151_/CLK _17996_/D vssd1 vssd1 vccd1 vccd1 _17996_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_215_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16947_ _18837_/Q _18801_/Q _16947_/S vssd1 vssd1 vccd1 vccd1 _16947_/X sky130_fd_sc_hd__mux2_1
XFILLER_133_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_226_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16878_ _17148_/A vssd1 vssd1 vccd1 vccd1 _16936_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_92_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_231_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18617_ _18620_/CLK _18617_/D vssd1 vssd1 vccd1 vccd1 _18617_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_168_1346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15829_ _15876_/A _15829_/B vssd1 vssd1 vccd1 vccd1 _15829_/Y sky130_fd_sc_hd__nand2_1
XFILLER_64_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09350_ _18437_/Q _18436_/Q _18435_/Q vssd1 vssd1 vccd1 vccd1 _09354_/A sky130_fd_sc_hd__or3_4
XFILLER_64_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18548_ _18548_/CLK _18548_/D vssd1 vssd1 vccd1 vccd1 _18548_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_209_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_178_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09281_ _18851_/Q _18850_/Q _18849_/Q vssd1 vssd1 vccd1 vccd1 _09282_/D sky130_fd_sc_hd__or3_2
X_18479_ _18482_/CLK _18479_/D vssd1 vssd1 vccd1 vccd1 _18479_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_127_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_220_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_1347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_1328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_142_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_5_28_0_wb_clk_i clkbuf_5_29_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_5_28_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_87_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08996_ _08997_/A vssd1 vssd1 vccd1 vccd1 _08996_/Y sky130_fd_sc_hd__inv_2
XFILLER_125_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_229_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_228_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_214_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_1266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_229_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09617_ _09617_/A _09617_/B vssd1 vssd1 vccd1 vccd1 _09618_/B sky130_fd_sc_hd__nand2_1
XFILLER_141_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_231_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09548_ _18103_/Q _10618_/A vssd1 vssd1 vccd1 vccd1 _09549_/B sky130_fd_sc_hd__xor2_1
XFILLER_70_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_231_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_180_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09479_ _09474_/Y _09467_/B _18138_/D vssd1 vssd1 vccd1 vccd1 _18144_/D sky130_fd_sc_hd__o21a_1
XFILLER_196_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_169_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_200_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_180_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11510_ _17871_/Q vssd1 vssd1 vccd1 vccd1 _11530_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_106_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12490_ _12490_/A _12495_/C _12490_/C vssd1 vssd1 vccd1 vccd1 _12491_/A sky130_fd_sc_hd__and3_1
XFILLER_106_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11441_ _11428_/Y _11440_/X _11828_/B vssd1 vssd1 vccd1 vccd1 _11441_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_109_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14160_ _18965_/Q _13493_/A _14030_/X _18980_/Q vssd1 vssd1 vccd1 vccd1 _14160_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_109_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11372_ _11582_/A _13446_/A vssd1 vssd1 vccd1 vccd1 _11374_/A sky130_fd_sc_hd__and2_1
XFILLER_50_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13111_ _13111_/A vssd1 vssd1 vccd1 vccd1 _18015_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_30_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10323_ _10321_/X _10322_/X _10598_/A vssd1 vssd1 vccd1 vccd1 _10323_/X sky130_fd_sc_hd__mux2_1
X_14091_ _18434_/Q _13848_/X _13858_/A _18425_/Q vssd1 vssd1 vccd1 vccd1 _14091_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_152_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_166_wb_clk_i clkbuf_5_10_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18085_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_3_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13042_ _17993_/Q _12783_/A _13025_/A _13041_/Y _13368_/B vssd1 vssd1 vccd1 vccd1
+ _13043_/B sky130_fd_sc_hd__a32o_1
XFILLER_112_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10254_ _10250_/X _11917_/A _10253_/X vssd1 vssd1 vccd1 vccd1 _10256_/A sky130_fd_sc_hd__a21oi_1
XFILLER_180_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_121_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17850_ _17891_/CLK _17850_/D vssd1 vssd1 vccd1 vccd1 _17850_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_65_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10185_ _10201_/A vssd1 vssd1 vccd1 vccd1 _10215_/A sky130_fd_sc_hd__buf_2
XFILLER_121_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16801_ _16803_/B _16798_/X _16799_/Y _16800_/X vssd1 vssd1 vccd1 vccd1 _18769_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_94_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_182_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17781_ _18110_/CLK _17781_/D vssd1 vssd1 vccd1 vccd1 _17781_/Q sky130_fd_sc_hd__dfxtp_2
X_14993_ _14995_/B _14991_/X _14992_/Y _14980_/X vssd1 vssd1 vccd1 vccd1 _18337_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_208_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16732_ _16755_/A _16732_/B vssd1 vssd1 vccd1 vccd1 _16732_/Y sky130_fd_sc_hd__nand2_1
XFILLER_219_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13944_ _18796_/Q _13529_/A _13725_/X _18772_/Q vssd1 vssd1 vccd1 vccd1 _13944_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_207_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13875_ _18481_/Q _13612_/X _13868_/X _13874_/X vssd1 vssd1 vccd1 vccd1 _13875_/X
+ sky130_fd_sc_hd__a211o_2
X_16663_ _16807_/A _16796_/C vssd1 vssd1 vccd1 vccd1 _16670_/B sky130_fd_sc_hd__nor2_2
XFILLER_74_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_228_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18402_ _18404_/CLK _18402_/D vssd1 vssd1 vccd1 vccd1 _18402_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_46_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_222_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15614_ _18483_/Q _15618_/B _15613_/X _15595_/X vssd1 vssd1 vccd1 vccd1 _18483_/D
+ sky130_fd_sc_hd__o211a_1
X_12826_ _12629_/A _12824_/Y _17957_/Q _12637_/B _12825_/X vssd1 vssd1 vccd1 vccd1
+ _12835_/A sky130_fd_sc_hd__o221ai_1
XFILLER_90_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16594_ _16599_/B _16592_/X _16593_/X _16581_/X vssd1 vssd1 vccd1 vccd1 _18717_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_37_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_188_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18333_ _18343_/CLK _18333_/D vssd1 vssd1 vccd1 vccd1 _18333_/Q sky130_fd_sc_hd__dfxtp_2
X_15545_ _18503_/Q _18467_/Q _15545_/S vssd1 vssd1 vccd1 vccd1 _15545_/X sky130_fd_sc_hd__mux2_1
X_12757_ _12920_/B _12920_/C vssd1 vssd1 vccd1 vccd1 _12757_/X sky130_fd_sc_hd__and2_1
XFILLER_15_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11708_ _11696_/C _11687_/Y _11703_/A vssd1 vssd1 vccd1 vccd1 _11708_/Y sky130_fd_sc_hd__a21oi_1
X_15476_ _15915_/A _15599_/C vssd1 vssd1 vccd1 vccd1 _15487_/B sky130_fd_sc_hd__nor2_2
X_18264_ _18266_/CLK _18264_/D vssd1 vssd1 vccd1 vccd1 _18264_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_124_1238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12688_ _12688_/A _12688_/B vssd1 vssd1 vccd1 vccd1 _12688_/Y sky130_fd_sc_hd__nand2_1
XFILLER_163_1298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_202_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14427_ _14422_/X _09499_/B _14423_/X vssd1 vssd1 vccd1 vccd1 _14427_/X sky130_fd_sc_hd__a21o_1
X_17215_ _17503_/A _17254_/B vssd1 vssd1 vccd1 vccd1 _17230_/B sky130_fd_sc_hd__nor2_2
XFILLER_175_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11639_ _11639_/A _11672_/A vssd1 vssd1 vccd1 vccd1 _11668_/A sky130_fd_sc_hd__nor2_1
XFILLER_204_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18195_ _18991_/CLK _18195_/D vssd1 vssd1 vccd1 vccd1 _18195_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_129_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14358_ _14203_/X _14355_/C _14355_/D _14357_/X vssd1 vssd1 vccd1 vccd1 _14358_/X
+ sky130_fd_sc_hd__o31a_1
X_17146_ _17435_/A _17202_/B vssd1 vssd1 vccd1 vccd1 _17156_/B sky130_fd_sc_hd__nor2_2
XFILLER_7_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13309_ _13309_/A _13309_/B _13309_/C vssd1 vssd1 vccd1 vccd1 _13310_/C sky130_fd_sc_hd__or3_1
X_17077_ _17080_/B _17074_/X _17075_/Y _17076_/X vssd1 vssd1 vccd1 vccd1 _18832_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_115_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14289_ _14289_/A _14307_/B vssd1 vssd1 vccd1 vccd1 _14289_/Y sky130_fd_sc_hd__nor2_1
XFILLER_170_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16028_ _16028_/A vssd1 vssd1 vccd1 vccd1 _16028_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_115_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_1334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17979_ _17990_/CLK _17979_/D vssd1 vssd1 vccd1 vccd1 _17979_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_211_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_226_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09402_ _09402_/A _09402_/B _10877_/A _09402_/D vssd1 vssd1 vccd1 vccd1 _09403_/C
+ sky130_fd_sc_hd__and4_1
XFILLER_129_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_213_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09333_ _18530_/Q _18529_/Q _18528_/Q vssd1 vssd1 vccd1 vccd1 _09337_/A sky130_fd_sc_hd__or3_4
XFILLER_34_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_221_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09264_ _18983_/Q _18982_/Q _18981_/Q vssd1 vssd1 vccd1 vccd1 _09265_/D sky130_fd_sc_hd__or3_2
XFILLER_139_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09195_ _18584_/Q _18583_/Q _18582_/Q vssd1 vssd1 vccd1 vccd1 _09198_/B sky130_fd_sc_hd__or3_4
XFILLER_14_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_140_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08979_ _08979_/A vssd1 vssd1 vccd1 vccd1 _08979_/Y sky130_fd_sc_hd__inv_2
XTAP_4825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19083__54 vssd1 vssd1 vccd1 vccd1 _19083__54/HI _19191_/A sky130_fd_sc_hd__conb_1
XTAP_4836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11990_ _12055_/C _12009_/C _11990_/C vssd1 vssd1 vccd1 vccd1 _13710_/B sky130_fd_sc_hd__and3b_2
XTAP_4869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_216_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10941_ _09392_/C _10069_/X _10940_/X _09360_/D _10944_/S vssd1 vssd1 vccd1 vccd1
+ _10941_/X sky130_fd_sc_hd__a221o_1
XFILLER_44_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_216_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13660_ _18981_/Q _13657_/X _13658_/X _13659_/X vssd1 vssd1 vccd1 vccd1 _13660_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_216_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_1238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10872_ _09408_/C _10644_/A _10871_/X _10693_/X vssd1 vssd1 vccd1 vccd1 _10872_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_71_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12611_ _12600_/A _12600_/B _12600_/C _12598_/B vssd1 vssd1 vccd1 vccd1 _12612_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_188_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_213_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13591_ _13869_/A vssd1 vssd1 vccd1 vccd1 _13591_/X sky130_fd_sc_hd__buf_6
XPHY_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_213_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15330_ _18453_/Q _18417_/Q _15334_/S vssd1 vssd1 vccd1 vccd1 _15330_/X sky130_fd_sc_hd__mux2_1
XPHY_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12542_ _12574_/B _12542_/B vssd1 vssd1 vccd1 vccd1 _12542_/Y sky130_fd_sc_hd__nand2_1
XFILLER_101_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_212_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15261_ _15263_/B _15259_/X _15260_/Y _15244_/X vssd1 vssd1 vccd1 vccd1 _18403_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_12_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12473_ _12473_/A vssd1 vssd1 vccd1 vccd1 _17906_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_138_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17000_ _16998_/B _16997_/X _16998_/Y _16999_/X vssd1 vssd1 vccd1 vccd1 _18812_/D
+ sky130_fd_sc_hd__o211a_1
X_14212_ _18213_/Q _18212_/Q _18206_/Q vssd1 vssd1 vccd1 vccd1 _14212_/X sky130_fd_sc_hd__or3b_1
X_11424_ _12329_/A _11419_/X _11645_/A _12323_/A _11423_/Y vssd1 vssd1 vccd1 vccd1
+ _11424_/X sky130_fd_sc_hd__o221a_1
XFILLER_6_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15192_ _15195_/B _15189_/X _15191_/Y _15187_/X vssd1 vssd1 vccd1 vccd1 _18385_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_184_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_1293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14143_ _18590_/Q _13575_/A _14026_/A _18581_/Q vssd1 vssd1 vccd1 vccd1 _14143_/X
+ sky130_fd_sc_hd__a22o_1
X_11355_ _11359_/B _17798_/Q _11403_/A vssd1 vssd1 vccd1 vccd1 _11453_/B sky130_fd_sc_hd__o21ai_2
XFILLER_67_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_1356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_1307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10306_ _09170_/A _09165_/D _09160_/D _09170_/C _10291_/A _10285_/S vssd1 vssd1 vccd1
+ vccd1 _10306_/X sky130_fd_sc_hd__mux4_1
X_14074_ _18716_/Q _13877_/X _13842_/A _18710_/Q vssd1 vssd1 vccd1 vccd1 _14074_/X
+ sky130_fd_sc_hd__a22o_1
X_18951_ _18953_/CLK _18951_/D vssd1 vssd1 vccd1 vccd1 _18951_/Q sky130_fd_sc_hd__dfxtp_1
X_11286_ _13447_/A _11404_/B vssd1 vssd1 vccd1 vccd1 _11286_/X sky130_fd_sc_hd__and2_1
X_17902_ _17911_/CLK _17902_/D vssd1 vssd1 vccd1 vccd1 _17902_/Q sky130_fd_sc_hd__dfxtp_1
X_13025_ _13025_/A vssd1 vssd1 vccd1 vccd1 _13025_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_112_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10237_ _10883_/A _09360_/C _09365_/A _09370_/B _10231_/X _10236_/X vssd1 vssd1 vccd1
+ vccd1 _10237_/X sky130_fd_sc_hd__mux4_2
X_18882_ _18907_/CLK _18882_/D vssd1 vssd1 vccd1 vccd1 _18882_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_6_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17833_ _18217_/CLK _17833_/D vssd1 vssd1 vccd1 vccd1 _17833_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_67_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10168_ _10162_/A _10168_/B vssd1 vssd1 vccd1 vccd1 _10169_/B sky130_fd_sc_hd__and2b_1
XFILLER_86_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17764_ _17764_/A _19026_/Q vssd1 vssd1 vccd1 vccd1 _17765_/A sky130_fd_sc_hd__and2_1
X_14976_ _14983_/B _14974_/X _14975_/X _14961_/X vssd1 vssd1 vccd1 vccd1 _18333_/D
+ sky130_fd_sc_hd__o211a_1
X_10099_ _10085_/S _10096_/X _10098_/X _10041_/A vssd1 vssd1 vccd1 vccd1 _10099_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_212_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_208_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_63_wb_clk_i clkbuf_5_20_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18710_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_16715_ _18783_/Q _18747_/Q _16715_/S vssd1 vssd1 vccd1 vccd1 _16715_/X sky130_fd_sc_hd__mux2_1
XFILLER_212_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13927_ _18235_/Q _13505_/A _13626_/A _18259_/Q vssd1 vssd1 vccd1 vccd1 _13927_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_223_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17695_ _17645_/X _17687_/Y _17552_/A _17688_/Y _18986_/Q vssd1 vssd1 vccd1 vccd1
+ _17696_/B sky130_fd_sc_hd__a32o_1
XFILLER_62_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_228_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16646_ _18767_/Q _18731_/Q _16657_/S vssd1 vssd1 vccd1 vccd1 _16646_/X sky130_fd_sc_hd__mux2_1
XFILLER_165_1327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13858_ _13858_/A vssd1 vssd1 vccd1 vccd1 _13858_/X sky130_fd_sc_hd__buf_4
XFILLER_62_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_223_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_204_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12809_ _12809_/A _17948_/Q vssd1 vssd1 vccd1 vccd1 _12809_/Y sky130_fd_sc_hd__nand2_1
X_16577_ _17037_/A _16652_/C vssd1 vssd1 vccd1 vccd1 _16589_/B sky130_fd_sc_hd__nor2_2
X_13789_ _18444_/Q _13759_/X _13780_/X _18435_/Q _13788_/X vssd1 vssd1 vccd1 vccd1
+ _13789_/X sky130_fd_sc_hd__a221o_4
XFILLER_96_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18316_ _18317_/CLK _18316_/D vssd1 vssd1 vccd1 vccd1 _18316_/Q sky130_fd_sc_hd__dfxtp_4
X_15528_ _16431_/A vssd1 vssd1 vccd1 vccd1 _16128_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_124_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18247_ _18809_/CLK _18247_/D vssd1 vssd1 vccd1 vccd1 _18247_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15459_ _15582_/A vssd1 vssd1 vccd1 vccd1 _15511_/A sky130_fd_sc_hd__buf_2
XFILLER_198_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18178_ _18178_/CLK _18178_/D vssd1 vssd1 vccd1 vccd1 _18178_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_191_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_1306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_1366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17129_ _17156_/A _17129_/B vssd1 vssd1 vccd1 vccd1 _17129_/Y sky130_fd_sc_hd__nand2_1
XFILLER_7_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09951_ _10600_/A vssd1 vssd1 vccd1 vccd1 _10391_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_116_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09882_ _09882_/A _09883_/B vssd1 vssd1 vccd1 vccd1 _09887_/B sky130_fd_sc_hd__xnor2_4
XFILLER_112_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_211_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_226_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_213_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09316_ _18470_/Q _18469_/Q _18468_/Q vssd1 vssd1 vccd1 vccd1 _09319_/B sky130_fd_sc_hd__or3_4
XFILLER_16_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_142_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09247_ _18881_/Q _18880_/Q _18879_/Q vssd1 vssd1 vccd1 vccd1 _10097_/A sky130_fd_sc_hd__or3_4
XFILLER_194_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09178_ _18620_/Q _18619_/Q _18618_/Q vssd1 vssd1 vccd1 vccd1 _09181_/B sky130_fd_sc_hd__or3_4
XFILLER_5_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_218_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11140_ _11498_/A vssd1 vssd1 vccd1 vccd1 _13485_/A sky130_fd_sc_hd__buf_2
XFILLER_1_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_6013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11071_ _11895_/A vssd1 vssd1 vccd1 vccd1 _11091_/S sky130_fd_sc_hd__clkbuf_2
XTAP_6046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10022_ _09126_/C _09131_/B _09136_/D _09131_/D _10955_/S _10065_/A vssd1 vssd1 vccd1
+ vccd1 _10022_/X sky130_fd_sc_hd__mux4_1
XFILLER_62_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14830_ _18333_/Q _18297_/Q _14830_/S vssd1 vssd1 vccd1 vccd1 _14830_/X sky130_fd_sc_hd__mux2_1
XFILLER_76_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14761_ _18316_/Q _18280_/Q _14787_/S vssd1 vssd1 vccd1 vccd1 _14761_/X sky130_fd_sc_hd__mux2_1
X_11973_ _11973_/A _11973_/B vssd1 vssd1 vccd1 vccd1 _13434_/A sky130_fd_sc_hd__and2_4
XTAP_4699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16500_ _16499_/B _16498_/X _16499_/Y _16496_/X vssd1 vssd1 vccd1 vccd1 _18695_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_3976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10924_ _10920_/X _10923_/X _12039_/A vssd1 vssd1 vccd1 vccd1 _10924_/X sky130_fd_sc_hd__mux2_1
X_13712_ _13637_/Y _13647_/X _13696_/X _13711_/X vssd1 vssd1 vccd1 vccd1 _13712_/X
+ sky130_fd_sc_hd__a211o_2
XFILLER_217_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14692_ _14778_/A vssd1 vssd1 vccd1 vccd1 _14692_/X sky130_fd_sc_hd__buf_4
XFILLER_45_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17480_ _17480_/A _17491_/B vssd1 vssd1 vccd1 vccd1 _17489_/B sky130_fd_sc_hd__nor2_2
XFILLER_186_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16431_ _16431_/A vssd1 vssd1 vccd1 vccd1 _17037_/A sky130_fd_sc_hd__buf_6
XFILLER_16_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10855_ _09370_/A _09360_/B _10870_/S vssd1 vssd1 vccd1 vccd1 _10855_/X sky130_fd_sc_hd__mux2_1
X_13643_ _18882_/Q _13642_/X _13861_/A _18906_/Q vssd1 vssd1 vccd1 vccd1 _13643_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_44_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_213_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19150_ _19150_/A _09036_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[20] sky130_fd_sc_hd__ebufn_8
XFILLER_198_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16362_ _16364_/B _16360_/X _16361_/Y _16354_/X vssd1 vssd1 vccd1 vccd1 _18661_/D
+ sky130_fd_sc_hd__o211a_1
X_13574_ _14081_/B vssd1 vssd1 vccd1 vccd1 _13575_/A sky130_fd_sc_hd__buf_6
XFILLER_160_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10786_ _10843_/C vssd1 vssd1 vccd1 vccd1 _10910_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_201_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18101_ _18130_/CLK _18101_/D vssd1 vssd1 vccd1 vccd1 _18101_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15313_ _15840_/A vssd1 vssd1 vccd1 vccd1 _15739_/A sky130_fd_sc_hd__clkbuf_2
X_12525_ _17919_/Q vssd1 vssd1 vccd1 vccd1 _12809_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_16293_ _18643_/Q _16294_/B _16292_/Y _16274_/X vssd1 vssd1 vccd1 vccd1 _18643_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_185_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_181_wb_clk_i clkbuf_5_8_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _19009_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_201_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_185_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18032_ _18035_/CLK _18032_/D vssd1 vssd1 vccd1 vccd1 _18032_/Q sky130_fd_sc_hd__dfxtp_1
X_15244_ _15283_/A vssd1 vssd1 vccd1 vccd1 _15244_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_12456_ _17904_/Q _12470_/B vssd1 vssd1 vccd1 vccd1 _12477_/B sky130_fd_sc_hd__xor2_2
Xclkbuf_leaf_110_wb_clk_i clkbuf_5_31_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18496_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_184_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11407_ _11498_/A _11541_/A vssd1 vssd1 vccd1 vccd1 _11617_/C sky130_fd_sc_hd__or2_1
XFILLER_193_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15175_ _15220_/A _15175_/B _15199_/C vssd1 vssd1 vccd1 vccd1 _15175_/X sky130_fd_sc_hd__or3_1
XFILLER_125_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12387_ _12387_/A vssd1 vssd1 vccd1 vccd1 _12490_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_207_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14126_ _18911_/Q _13617_/X _14123_/X _14125_/X vssd1 vssd1 vccd1 vccd1 _14126_/X
+ sky130_fd_sc_hd__a211o_1
X_11338_ _11338_/A vssd1 vssd1 vccd1 vccd1 _11339_/B sky130_fd_sc_hd__clkbuf_4
Xclkbuf_4_9_0_wb_clk_i clkbuf_4_9_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_4_9_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_45_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14057_ _18518_/Q _13612_/A _13576_/A _18509_/Q _14056_/X vssd1 vssd1 vccd1 vccd1
+ _14057_/X sky130_fd_sc_hd__a221o_1
X_18934_ _18936_/CLK _18934_/D vssd1 vssd1 vccd1 vccd1 _18934_/Q sky130_fd_sc_hd__dfxtp_4
X_11269_ _17791_/Q _17792_/Q vssd1 vssd1 vccd1 vccd1 _11926_/B sky130_fd_sc_hd__or2_1
XFILLER_45_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13008_ _13007_/B _13006_/X _13007_/Y _12964_/X vssd1 vssd1 vccd1 vccd1 _17981_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_80_1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_1364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18865_ _18865_/CLK _18865_/D vssd1 vssd1 vccd1 vccd1 _18865_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_228_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17816_ _17817_/CLK _17816_/D vssd1 vssd1 vccd1 vccd1 _17816_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_11_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18796_ _18812_/CLK _18796_/D vssd1 vssd1 vccd1 vccd1 _18796_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_67_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17747_ _17747_/A vssd1 vssd1 vccd1 vccd1 _17756_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_36_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14959_ _18365_/Q _18329_/Q _14974_/S vssd1 vssd1 vccd1 vccd1 _14959_/X sky130_fd_sc_hd__mux2_1
XFILLER_47_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17678_ _17681_/A _17678_/B vssd1 vssd1 vccd1 vccd1 _17679_/A sky130_fd_sc_hd__and2_1
XINSDIODE2_220 _13834_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINSDIODE2_231 _15255_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XINSDIODE2_242 _18349_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16629_ _16634_/B _16626_/X _16628_/X _16619_/X vssd1 vssd1 vccd1 vccd1 _18726_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_165_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XINSDIODE2_253 _14457_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_196_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_264 _14436_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09101_ _18803_/Q _18802_/Q _18801_/Q vssd1 vssd1 vccd1 vccd1 _09103_/C sky130_fd_sc_hd__or3_4
XFILLER_31_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09032_ _09034_/A vssd1 vssd1 vccd1 vccd1 _09032_/Y sky130_fd_sc_hd__inv_2
XFILLER_108_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09934_ _10292_/S vssd1 vssd1 vccd1 vccd1 _10316_/S sky130_fd_sc_hd__buf_4
XFILLER_58_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09865_ _18124_/Q _09867_/B _09867_/A vssd1 vssd1 vccd1 vccd1 _09875_/A sky130_fd_sc_hd__a21bo_1
XFILLER_98_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_213_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19053__24 vssd1 vssd1 vccd1 vccd1 _19053__24/HI _19147_/A sky130_fd_sc_hd__conb_1
X_09796_ _09816_/B _09816_/C _09816_/A vssd1 vssd1 vccd1 vccd1 _09817_/B sky130_fd_sc_hd__a21oi_1
XTAP_3206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10640_ _10640_/A _10656_/B vssd1 vssd1 vccd1 vccd1 _10716_/A sky130_fd_sc_hd__xnor2_4
XFILLER_195_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10571_ _10090_/S _10567_/X _10570_/X _10893_/S vssd1 vssd1 vccd1 vccd1 _10571_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_107_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_220_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12310_ _11323_/X _12292_/B _11346_/A vssd1 vssd1 vccd1 vccd1 _12311_/C sky130_fd_sc_hd__a21o_1
XFILLER_107_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13290_ _19026_/Q _19025_/Q _18011_/Q _18010_/Q vssd1 vssd1 vccd1 vccd1 _13291_/D
+ sky130_fd_sc_hd__or4_1
XFILLER_213_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12241_ _17859_/Q _17858_/Q _12223_/X vssd1 vssd1 vccd1 vccd1 _12269_/B sky130_fd_sc_hd__o21a_2
XFILLER_108_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12172_ _17845_/Q _12172_/B vssd1 vssd1 vccd1 vccd1 _12172_/X sky130_fd_sc_hd__and2_1
XFILLER_122_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_218_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11123_ _11123_/A vssd1 vssd1 vccd1 vccd1 _17798_/D sky130_fd_sc_hd__clkbuf_1
X_16980_ _14354_/X _16975_/X _16978_/X _16979_/Y _14618_/X vssd1 vssd1 vccd1 vccd1
+ _18807_/D sky130_fd_sc_hd__o311a_1
XFILLER_104_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15931_ _15931_/A _15993_/B vssd1 vssd1 vccd1 vccd1 _15942_/B sky130_fd_sc_hd__nor2_2
XTAP_5120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11054_ _11333_/A _11215_/B _12272_/A vssd1 vssd1 vccd1 vccd1 _11055_/A sky130_fd_sc_hd__mux2_1
XFILLER_107_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10005_ _09109_/A _10003_/S _10004_/X _09987_/X vssd1 vssd1 vccd1 vccd1 _10005_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_209_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18650_ _18650_/CLK _18650_/D vssd1 vssd1 vccd1 vccd1 _18650_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_5164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15862_ _15865_/B _15859_/X _15860_/Y _15861_/X vssd1 vssd1 vccd1 vccd1 _18544_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_190_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17601_ _17601_/A vssd1 vssd1 vccd1 vccd1 _18962_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_190_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14813_ _18329_/Q _18293_/Q _14830_/S vssd1 vssd1 vccd1 vccd1 _14813_/X sky130_fd_sc_hd__mux2_1
X_18581_ _18593_/CLK _18581_/D vssd1 vssd1 vccd1 vccd1 _18581_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_4474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15793_ _15863_/A vssd1 vssd1 vccd1 vccd1 _15809_/S sky130_fd_sc_hd__buf_2
XTAP_4485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_229_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17532_ _17534_/B _17530_/X _17531_/Y _17517_/X vssd1 vssd1 vccd1 vccd1 _18946_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_3773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14744_ _15184_/A _14790_/B vssd1 vssd1 vccd1 vccd1 _14753_/B sky130_fd_sc_hd__nor2_2
XFILLER_17_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11956_ _12049_/A _11960_/C _11939_/X _11944_/X vssd1 vssd1 vccd1 vccd1 _11957_/B
+ sky130_fd_sc_hd__o211a_4
XTAP_3795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_229_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_205_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17463_ _18964_/Q _18928_/Q _17467_/S vssd1 vssd1 vccd1 vccd1 _17463_/X sky130_fd_sc_hd__mux2_1
X_10907_ _09376_/A _09386_/B _09381_/A _09376_/D _14206_/A _10852_/X vssd1 vssd1 vccd1
+ vccd1 _10907_/X sky130_fd_sc_hd__mux4_1
X_14675_ _17575_/A vssd1 vssd1 vccd1 vccd1 _14928_/A sky130_fd_sc_hd__clkbuf_2
X_11887_ _12207_/A _11887_/B vssd1 vssd1 vccd1 vccd1 _17835_/D sky130_fd_sc_hd__nor2_1
XFILLER_44_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19202_ _19202_/A _08987_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[2] sky130_fd_sc_hd__ebufn_8
X_16414_ _16447_/A _16417_/B vssd1 vssd1 vccd1 vccd1 _16414_/Y sky130_fd_sc_hd__nand2_1
XFILLER_189_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13626_ _13626_/A vssd1 vssd1 vccd1 vccd1 _13703_/A sky130_fd_sc_hd__buf_4
XFILLER_20_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10838_ _10838_/A _10838_/B _10838_/C vssd1 vssd1 vccd1 vccd1 _10838_/X sky130_fd_sc_hd__or3_1
X_17394_ _18947_/Q _18911_/Q _17406_/S vssd1 vssd1 vccd1 vccd1 _17394_/X sky130_fd_sc_hd__mux2_1
XFILLER_186_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19133_ _19133_/A _09051_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[3] sky130_fd_sc_hd__ebufn_8
XFILLER_201_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16345_ _18693_/Q _18657_/Q _16345_/S vssd1 vssd1 vccd1 vccd1 _16345_/X sky130_fd_sc_hd__mux2_1
XFILLER_201_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13557_ _13557_/A _13557_/B vssd1 vssd1 vccd1 vccd1 _13583_/A sky130_fd_sc_hd__nor2_8
X_10769_ _10838_/A _10671_/B _10768_/Y _12101_/A _10843_/B vssd1 vssd1 vccd1 vccd1
+ _10773_/B sky130_fd_sc_hd__a311o_1
XFILLER_121_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12508_ _12521_/A _12528_/C vssd1 vssd1 vccd1 vccd1 _12514_/A sky130_fd_sc_hd__or2_1
X_16276_ _16327_/A vssd1 vssd1 vccd1 vccd1 _16304_/S sky130_fd_sc_hd__clkbuf_2
X_13488_ _13652_/A vssd1 vssd1 vccd1 vccd1 _13489_/A sky130_fd_sc_hd__buf_6
XFILLER_145_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18015_ _19004_/CLK _18015_/D vssd1 vssd1 vccd1 vccd1 _18015_/Q sky130_fd_sc_hd__dfxtp_1
X_15227_ _15239_/A _15227_/B vssd1 vssd1 vccd1 vccd1 _15227_/Y sky130_fd_sc_hd__nand2_1
X_12439_ _12439_/A _12439_/B _12439_/C _12439_/D vssd1 vssd1 vccd1 vccd1 _12440_/B
+ sky130_fd_sc_hd__nand4_1
XFILLER_201_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15158_ _18147_/Q _15772_/B vssd1 vssd1 vccd1 vccd1 _15270_/A sky130_fd_sc_hd__nand2_4
XFILLER_141_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14109_ _18779_/Q _13577_/X _14105_/X _14108_/X vssd1 vssd1 vccd1 vccd1 _14109_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_99_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15089_ _15094_/B _15087_/X _15088_/X _15083_/X vssd1 vssd1 vccd1 vccd1 _18360_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_99_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18917_ _18931_/CLK _18917_/D vssd1 vssd1 vccd1 vccd1 _18917_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_132_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09650_ _09649_/B _09704_/A _09649_/A vssd1 vssd1 vccd1 vccd1 _09679_/A sky130_fd_sc_hd__o21a_1
XFILLER_227_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18848_ _18866_/CLK _18848_/D vssd1 vssd1 vccd1 vccd1 _18848_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_110_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_216_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09581_ _09565_/A _09565_/B _09580_/X vssd1 vssd1 vccd1 vccd1 _09600_/C sky130_fd_sc_hd__a21o_1
X_18779_ _18786_/CLK _18779_/D vssd1 vssd1 vccd1 vccd1 _18779_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_94_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_223_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_211_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_1290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_136_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_192_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09015_ _09016_/A vssd1 vssd1 vccd1 vccd1 _09015_/Y sky130_fd_sc_hd__inv_4
XFILLER_163_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_219_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_117_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09917_ _09895_/X _09906_/X _09914_/X _09916_/X vssd1 vssd1 vccd1 vccd1 _09932_/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_104_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09848_ _17781_/Q _10193_/B vssd1 vssd1 vccd1 vccd1 _09853_/A sky130_fd_sc_hd__xnor2_2
XFILLER_24_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09779_ _10213_/A _09780_/B vssd1 vssd1 vccd1 vccd1 _09779_/X sky130_fd_sc_hd__or2_1
XTAP_3047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11810_ _11779_/X _11809_/X _11820_/A vssd1 vssd1 vccd1 vccd1 _11810_/X sky130_fd_sc_hd__o21a_1
XTAP_2324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12790_ _17944_/Q _13066_/C _12789_/X _12510_/X vssd1 vssd1 vccd1 vccd1 _17944_/D
+ sky130_fd_sc_hd__a211o_1
XTAP_2335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11741_ _11404_/B _11593_/A _11720_/A vssd1 vssd1 vccd1 vccd1 _11741_/X sky130_fd_sc_hd__a21o_1
XTAP_2368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_230_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11672_ _11672_/A _11672_/B vssd1 vssd1 vccd1 vccd1 _11673_/B sky130_fd_sc_hd__nand2_1
XTAP_1678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14460_ _14279_/A _17709_/B _14459_/Y vssd1 vssd1 vccd1 vccd1 _18206_/D sky130_fd_sc_hd__a21oi_1
XFILLER_144_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_1330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13411_ _13411_/A _13411_/B _13411_/C _13411_/D vssd1 vssd1 vccd1 vccd1 _13412_/B
+ sky130_fd_sc_hd__nor4_2
X_10623_ _10623_/A vssd1 vssd1 vccd1 vccd1 _12966_/A sky130_fd_sc_hd__buf_6
X_14391_ _18190_/Q _18189_/Q vssd1 vssd1 vccd1 vccd1 _14391_/Y sky130_fd_sc_hd__nor2_1
XFILLER_128_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16130_ _16130_/A _16132_/B vssd1 vssd1 vccd1 vccd1 _16130_/Y sky130_fd_sc_hd__nand2_1
XFILLER_155_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13342_ _13398_/A vssd1 vssd1 vccd1 vccd1 _13342_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_183_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10554_ _09181_/B _09176_/C _09186_/D _09176_/A _10494_/A _10522_/A vssd1 vssd1 vccd1
+ vccd1 _10555_/B sky130_fd_sc_hd__mux4_1
XFILLER_10_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_182_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16061_ _18591_/Q _16064_/B _16060_/X _16048_/X vssd1 vssd1 vccd1 vccd1 _18591_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_183_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13273_ _12987_/A _12747_/B _13272_/X _11896_/X _12748_/B vssd1 vssd1 vccd1 vccd1
+ _18089_/D sky130_fd_sc_hd__o2111a_1
XFILLER_170_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10485_ _09114_/A _09109_/A _09119_/B _10728_/A _10484_/X _10231_/X vssd1 vssd1 vccd1
+ vccd1 _10485_/X sky130_fd_sc_hd__mux4_2
XFILLER_120_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15012_ _15061_/A _15012_/B vssd1 vssd1 vccd1 vccd1 _15012_/Y sky130_fd_sc_hd__nand2_1
X_12224_ _12224_/A vssd1 vssd1 vccd1 vccd1 _12708_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_120_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_159_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12155_ _17842_/Q _12171_/B _12175_/B _11863_/X vssd1 vssd1 vccd1 vccd1 _17842_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_78_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11106_ _11720_/B _17806_/Q _11113_/S vssd1 vssd1 vccd1 vccd1 _11107_/A sky130_fd_sc_hd__mux2_1
XFILLER_111_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16963_ _17015_/A _17538_/B _16963_/C vssd1 vssd1 vccd1 vccd1 _16963_/X sky130_fd_sc_hd__or3_1
X_12086_ _14317_/B _12133_/B vssd1 vssd1 vccd1 vccd1 _12086_/X sky130_fd_sc_hd__or2_1
XFILLER_110_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_231_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18702_ _18708_/CLK _18702_/D vssd1 vssd1 vccd1 vccd1 _18702_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_204_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15914_ _18557_/Q _15913_/B _15913_/Y _15901_/X vssd1 vssd1 vccd1 vccd1 _18557_/D
+ sky130_fd_sc_hd__o211a_1
X_11037_ _17997_/Q _17996_/Q _11037_/C vssd1 vssd1 vccd1 vccd1 _13370_/B sky130_fd_sc_hd__and3_4
XFILLER_209_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16894_ _16903_/B _16888_/X _16890_/X _16893_/X vssd1 vssd1 vccd1 vccd1 _18789_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_37_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_231_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18633_ _18633_/CLK _18633_/D vssd1 vssd1 vccd1 vccd1 _18633_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_49_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_225_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15845_ _15863_/A vssd1 vssd1 vccd1 vccd1 _15859_/S sky130_fd_sc_hd__clkbuf_2
XTAP_4260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18564_ _18571_/CLK _18564_/D vssd1 vssd1 vccd1 vccd1 _18564_/Q sky130_fd_sc_hd__dfxtp_4
X_15776_ _15799_/A _15921_/B _15811_/C vssd1 vssd1 vccd1 vccd1 _15776_/X sky130_fd_sc_hd__or3_1
XTAP_3570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_220_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12988_ _12747_/B _12987_/Y _12927_/Y vssd1 vssd1 vccd1 vccd1 _12989_/A sky130_fd_sc_hd__a21bo_1
XFILLER_92_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17515_ _18978_/Q _18942_/Q _17515_/S vssd1 vssd1 vccd1 vccd1 _17515_/X sky130_fd_sc_hd__mux2_1
XFILLER_166_1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14727_ _14729_/B _14725_/X _14726_/Y _14716_/X vssd1 vssd1 vccd1 vccd1 _18271_/D
+ sky130_fd_sc_hd__o211a_1
X_18495_ _18497_/CLK _18495_/D vssd1 vssd1 vccd1 vccd1 _18495_/Q sky130_fd_sc_hd__dfxtp_2
X_11939_ _11929_/X _12007_/B _11937_/X _12015_/A vssd1 vssd1 vccd1 vccd1 _11939_/X
+ sky130_fd_sc_hd__o31a_2
XFILLER_162_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17446_ _17446_/A _17491_/B vssd1 vssd1 vccd1 vccd1 _17456_/B sky130_fd_sc_hd__nor2_1
XFILLER_220_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14658_ _14683_/A _14658_/B vssd1 vssd1 vccd1 vccd1 _14658_/Y sky130_fd_sc_hd__nand2_1
XFILLER_32_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_221_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13609_ _18807_/Q _13539_/X _13603_/X _13608_/X vssd1 vssd1 vccd1 vccd1 _13609_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_220_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17377_ _17383_/B _17375_/X _17376_/X _17361_/X vssd1 vssd1 vccd1 vccd1 _18906_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_158_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14589_ _14606_/A _14589_/B vssd1 vssd1 vccd1 vccd1 _14589_/Y sky130_fd_sc_hd__nand2_1
XFILLER_229_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16328_ _18689_/Q _18653_/Q _16345_/S vssd1 vssd1 vccd1 vccd1 _16328_/X sky130_fd_sc_hd__mux2_1
XFILLER_192_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_229_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_185_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16259_ _18672_/Q _18636_/Q _16271_/S vssd1 vssd1 vccd1 vccd1 _16259_/X sky130_fd_sc_hd__mux2_1
XFILLER_145_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_5_18_0_wb_clk_i clkbuf_4_9_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_5_18_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_88_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_8 _09119_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_228_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_214_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09702_ _09987_/A vssd1 vssd1 vccd1 vccd1 _09703_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_114_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_228_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_228_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_214_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_216_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09633_ _18098_/Q _12946_/A vssd1 vssd1 vccd1 vccd1 _09645_/B sky130_fd_sc_hd__xor2_1
XFILLER_215_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09564_ _18103_/Q _17980_/Q vssd1 vssd1 vccd1 vccd1 _09565_/B sky130_fd_sc_hd__xor2_1
Xclkbuf_leaf_213_wb_clk_i clkbuf_5_9_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17824_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_215_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09495_ _18192_/Q _09495_/B vssd1 vssd1 vccd1 vccd1 _14409_/B sky130_fd_sc_hd__or2_1
XFILLER_51_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_224_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_208_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_1268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_180_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_223_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_212_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_221_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_221_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_180_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10270_ _10270_/A _10270_/B _10270_/C vssd1 vssd1 vccd1 vccd1 _10271_/C sky130_fd_sc_hd__and3_1
XFILLER_191_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_219_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13960_ _18658_/Q _13615_/A _13958_/X _13959_/X vssd1 vssd1 vccd1 vccd1 _13960_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_59_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_219_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12911_ _12913_/A _12913_/C _12874_/X vssd1 vssd1 vccd1 vccd1 _12911_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_86_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_207_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13891_ _18613_/Q _13559_/A _13490_/A _18604_/Q vssd1 vssd1 vccd1 vccd1 _13891_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_24_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15630_ _15630_/A _15633_/B vssd1 vssd1 vccd1 vccd1 _15630_/Y sky130_fd_sc_hd__nand2_1
XFILLER_189_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12842_ _17945_/Q _17946_/Q vssd1 vssd1 vccd1 vccd1 _12846_/B sky130_fd_sc_hd__nand2_1
XTAP_2121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15561_ _18507_/Q _18471_/Q _15565_/S vssd1 vssd1 vccd1 vccd1 _15561_/X sky130_fd_sc_hd__mux2_1
XFILLER_27_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12773_ _13269_/B _12924_/B _12771_/Y _12772_/Y _12346_/A vssd1 vssd1 vccd1 vccd1
+ _17941_/D sky130_fd_sc_hd__a311oi_1
XTAP_1431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_215_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17300_ _17303_/B _17298_/X _17299_/Y _17283_/X vssd1 vssd1 vccd1 vccd1 _18886_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_9_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14512_ _14515_/B _14513_/B vssd1 vssd1 vccd1 vccd1 _14512_/Y sky130_fd_sc_hd__nor2_1
XTAP_2198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18280_ _18290_/CLK _18280_/D vssd1 vssd1 vccd1 vccd1 _18280_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_15_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11724_ _17912_/Q vssd1 vssd1 vccd1 vccd1 _11737_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_15492_ _15492_/A _15935_/B _15515_/C vssd1 vssd1 vccd1 vccd1 _15492_/X sky130_fd_sc_hd__or3_1
XTAP_1475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17231_ _17230_/B _17227_/X _17230_/Y _17219_/X vssd1 vssd1 vccd1 vccd1 _18869_/D
+ sky130_fd_sc_hd__o211a_1
X_11655_ _11795_/A _11655_/B _11655_/C _11442_/B vssd1 vssd1 vccd1 vccd1 _11665_/B
+ sky130_fd_sc_hd__or4b_2
X_14443_ _18201_/Q _14442_/X _14428_/X _14445_/B vssd1 vssd1 vccd1 vccd1 _14444_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_187_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_88_wb_clk_i _18144_/CLK vssd1 vssd1 vccd1 vccd1 _18658_/CLK sky130_fd_sc_hd__clkbuf_16
X_10606_ _10618_/A vssd1 vssd1 vccd1 vccd1 _13000_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_80_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17162_ _17169_/B _17159_/X _17160_/X _17161_/X vssd1 vssd1 vccd1 vccd1 _18852_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_128_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11586_ _11586_/A _11748_/B _11586_/C _11586_/D vssd1 vssd1 vccd1 vccd1 _11586_/X
+ sky130_fd_sc_hd__or4_1
X_14374_ _14370_/Y _14371_/X _14373_/X _14185_/A vssd1 vssd1 vccd1 vccd1 _18186_/D
+ sky130_fd_sc_hd__o31a_1
XFILLER_80_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_196_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16113_ _18639_/Q _18603_/Q _16113_/S vssd1 vssd1 vccd1 vccd1 _16113_/X sky130_fd_sc_hd__mux2_1
X_10537_ _09386_/B _09376_/D _09376_/A _09381_/A _10522_/A _10429_/X vssd1 vssd1 vccd1
+ vccd1 _10538_/B sky130_fd_sc_hd__mux4_2
XFILLER_116_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13325_ _18092_/Q _13313_/X _13324_/Y _13074_/X vssd1 vssd1 vccd1 vccd1 _18092_/D
+ sky130_fd_sc_hd__o211a_1
Xclkbuf_leaf_17_wb_clk_i clkbuf_5_5_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18866_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_183_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17093_ _17526_/A _17107_/B vssd1 vssd1 vccd1 vccd1 _17105_/B sky130_fd_sc_hd__nor2_2
XFILLER_183_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_1207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16044_ _16051_/B _16042_/X _16043_/X _16028_/X vssd1 vssd1 vccd1 vccd1 _18588_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_109_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_143_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13256_ _13256_/A vssd1 vssd1 vccd1 vccd1 _18081_/D sky130_fd_sc_hd__clkbuf_1
X_10468_ _10270_/A _10467_/X _10936_/S vssd1 vssd1 vccd1 vccd1 _10468_/X sky130_fd_sc_hd__a21bo_1
XFILLER_108_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19089__60 vssd1 vssd1 vccd1 vccd1 _19089__60/HI _19197_/A sky130_fd_sc_hd__conb_1
XFILLER_124_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12207_ _12207_/A _12207_/B vssd1 vssd1 vccd1 vccd1 _17851_/D sky130_fd_sc_hd__nor2_1
X_13187_ _13187_/A vssd1 vssd1 vccd1 vccd1 _18050_/D sky130_fd_sc_hd__clkbuf_1
X_10399_ _12131_/A _10399_/B _12133_/A vssd1 vssd1 vccd1 vccd1 _10399_/X sky130_fd_sc_hd__or3b_1
XFILLER_215_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12138_ _17942_/Q _18166_/Q _12144_/S vssd1 vssd1 vccd1 vccd1 _12139_/A sky130_fd_sc_hd__mux2_2
XFILLER_96_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17995_ _18061_/CLK _17995_/D vssd1 vssd1 vccd1 vccd1 _17995_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16946_ _17526_/A _16960_/B vssd1 vssd1 vccd1 vccd1 _16957_/B sky130_fd_sc_hd__nor2_2
X_12069_ _12069_/A _12069_/B _12069_/C _12069_/D vssd1 vssd1 vccd1 vccd1 _12069_/X
+ sky130_fd_sc_hd__or4_1
XFILLER_96_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16877_ _18182_/Q vssd1 vssd1 vccd1 vccd1 _17148_/A sky130_fd_sc_hd__buf_2
XFILLER_49_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_226_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_1208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18616_ _18620_/CLK _18616_/D vssd1 vssd1 vccd1 vccd1 _18616_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_92_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15828_ _15889_/A vssd1 vssd1 vccd1 vccd1 _15876_/A sky130_fd_sc_hd__buf_2
XTAP_4090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_225_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_231_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_1358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_213_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18547_ _18548_/CLK _18547_/D vssd1 vssd1 vccd1 vccd1 _18547_/Q sky130_fd_sc_hd__dfxtp_1
X_15759_ _16055_/A _15894_/C vssd1 vssd1 vccd1 vccd1 _15769_/B sky130_fd_sc_hd__nor2_2
XFILLER_33_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09280_ _18869_/Q _18868_/Q _18867_/Q vssd1 vssd1 vccd1 vccd1 _09282_/C sky130_fd_sc_hd__or3_4
XFILLER_205_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18478_ _18482_/CLK _18478_/D vssd1 vssd1 vccd1 vccd1 _18478_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_221_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_220_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17429_ _17432_/B _17427_/X _17428_/Y _17421_/X vssd1 vssd1 vccd1 vccd1 _18919_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_193_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_216_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08995_ _08997_/A vssd1 vssd1 vccd1 vccd1 _08995_/Y sky130_fd_sc_hd__inv_2
XFILLER_134_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_1340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_214_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_205_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_217_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09616_ _09822_/A _09617_/B _09617_/A vssd1 vssd1 vccd1 vccd1 _09668_/A sky130_fd_sc_hd__a21bo_4
XFILLER_44_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_231_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_225_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09547_ _17979_/Q vssd1 vssd1 vccd1 vccd1 _10618_/A sky130_fd_sc_hd__buf_2
XFILLER_93_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09478_ _18146_/D _09457_/B _18142_/D vssd1 vssd1 vccd1 vccd1 _18143_/D sky130_fd_sc_hd__o21a_1
XFILLER_145_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_4_11_0_wb_clk_i clkbuf_3_5_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_5_23_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_157_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_221_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11440_ _11423_/A _12323_/A _12323_/B _11431_/B _11431_/A vssd1 vssd1 vccd1 vccd1
+ _11440_/X sky130_fd_sc_hd__a311o_1
XFILLER_7_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_221_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11371_ _11347_/X _11371_/B vssd1 vssd1 vccd1 vccd1 _11371_/X sky130_fd_sc_hd__and2b_1
XFILLER_109_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13110_ _13118_/A _18016_/Q vssd1 vssd1 vccd1 vccd1 _13111_/A sky130_fd_sc_hd__and2_1
XFILLER_50_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10322_ _09287_/A _09287_/D _09282_/D _09282_/B _09937_/A _10316_/S vssd1 vssd1 vccd1
+ vccd1 _10322_/X sky130_fd_sc_hd__mux4_1
X_14090_ _18431_/Q _13525_/X _14017_/X _18419_/Q vssd1 vssd1 vccd1 vccd1 _14090_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_166_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13041_ _13041_/A _13041_/B vssd1 vssd1 vccd1 vccd1 _13041_/Y sky130_fd_sc_hd__nor2_2
XFILLER_69_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10253_ _10253_/A _13348_/A _10829_/A vssd1 vssd1 vccd1 vccd1 _10253_/X sky130_fd_sc_hd__and3_1
XFILLER_133_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10184_ _18128_/Q vssd1 vssd1 vccd1 vccd1 _10201_/A sky130_fd_sc_hd__inv_2
XFILLER_191_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16800_ _16871_/A vssd1 vssd1 vccd1 vccd1 _16800_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_78_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17780_ _18191_/CLK _17780_/D vssd1 vssd1 vccd1 vccd1 _17780_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_135_wb_clk_i clkbuf_5_27_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18343_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_14992_ _14992_/A _14995_/B vssd1 vssd1 vccd1 vccd1 _14992_/Y sky130_fd_sc_hd__nand2_1
XFILLER_59_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16731_ _18751_/Q _16732_/B _16730_/Y _16724_/X vssd1 vssd1 vccd1 vccd1 _18751_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_115_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13943_ _18775_/Q _13719_/X _13752_/X _18781_/Q vssd1 vssd1 vccd1 vccd1 _13943_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_19_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16662_ _16727_/A vssd1 vssd1 vccd1 vccd1 _16796_/C sky130_fd_sc_hd__buf_2
X_13874_ _18466_/Q _13525_/A _13621_/X _18469_/Q _13873_/X vssd1 vssd1 vccd1 vccd1
+ _13874_/X sky130_fd_sc_hd__a221o_1
XFILLER_46_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18401_ _18432_/CLK _18401_/D vssd1 vssd1 vccd1 vccd1 _18401_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_90_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15613_ _15613_/A _15909_/B _15666_/C vssd1 vssd1 vccd1 vccd1 _15613_/X sky130_fd_sc_hd__or3_1
XFILLER_61_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12825_ _12662_/B _12815_/Y _17963_/Q _12662_/A vssd1 vssd1 vccd1 vccd1 _12825_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_216_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16593_ _16615_/A _16736_/B _16628_/C vssd1 vssd1 vccd1 vccd1 _16593_/X sky130_fd_sc_hd__or3_1
XFILLER_201_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18332_ _18343_/CLK _18332_/D vssd1 vssd1 vccd1 vccd1 _18332_/Q sky130_fd_sc_hd__dfxtp_2
X_15544_ _15546_/B _15542_/X _15543_/Y _15536_/X vssd1 vssd1 vccd1 vccd1 _18466_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_163_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12756_ _18021_/Q _18020_/Q _18023_/Q _18022_/Q vssd1 vssd1 vccd1 vccd1 _12920_/C
+ sky130_fd_sc_hd__and4_1
XFILLER_30_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18263_ _18263_/CLK _18263_/D vssd1 vssd1 vccd1 vccd1 _18263_/Q sky130_fd_sc_hd__dfxtp_1
X_11707_ _11704_/A _11706_/Y _11685_/X vssd1 vssd1 vccd1 vccd1 _11707_/Y sky130_fd_sc_hd__a21oi_1
XTAP_1294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15475_ _18449_/Q _15473_/B _15473_/Y _15474_/X vssd1 vssd1 vccd1 vccd1 _18449_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_175_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12687_ _12672_/A _12672_/B _12679_/A _12686_/X vssd1 vssd1 vccd1 vccd1 _12688_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_204_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17214_ _17213_/B _17212_/X _17213_/Y _17197_/X vssd1 vssd1 vccd1 vccd1 _18866_/D
+ sky130_fd_sc_hd__o211a_1
X_14426_ _14452_/A _14426_/B vssd1 vssd1 vccd1 vccd1 _18196_/D sky130_fd_sc_hd__nor2_1
XFILLER_198_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11638_ _17862_/Q _19035_/Q vssd1 vssd1 vccd1 vccd1 _11672_/A sky130_fd_sc_hd__or2b_1
X_18194_ _18991_/CLK _18194_/D vssd1 vssd1 vccd1 vccd1 _18194_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_200_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_204_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17145_ _17184_/A vssd1 vssd1 vccd1 vccd1 _17202_/B sky130_fd_sc_hd__buf_2
XFILLER_7_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14357_ _18183_/Q vssd1 vssd1 vccd1 vccd1 _14357_/X sky130_fd_sc_hd__buf_4
XFILLER_200_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11569_ _17867_/Q _11569_/B vssd1 vssd1 vccd1 vccd1 _11570_/B sky130_fd_sc_hd__and2_1
XFILLER_155_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13308_ _18085_/Q _18084_/Q _18087_/Q _18086_/Q vssd1 vssd1 vccd1 vccd1 _13309_/C
+ sky130_fd_sc_hd__or4_1
XFILLER_143_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17076_ _17096_/A vssd1 vssd1 vccd1 vccd1 _17076_/X sky130_fd_sc_hd__clkbuf_2
X_14288_ _18996_/Q _14204_/B vssd1 vssd1 vccd1 vccd1 _14307_/B sky130_fd_sc_hd__or2b_1
XFILLER_100_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16027_ _16064_/A _16027_/B vssd1 vssd1 vccd1 vccd1 _16027_/Y sky130_fd_sc_hd__nand2_1
X_13239_ _13239_/A vssd1 vssd1 vccd1 vccd1 _18073_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_41_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_1215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17978_ _17990_/CLK _17978_/D vssd1 vssd1 vccd1 vccd1 _17978_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_69_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16929_ _18833_/Q _18797_/Q _16947_/S vssd1 vssd1 vccd1 vccd1 _16929_/X sky130_fd_sc_hd__mux2_1
XFILLER_211_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_226_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09401_ _18368_/Q _18367_/Q _18366_/Q vssd1 vssd1 vccd1 vccd1 _09402_/D sky130_fd_sc_hd__or3_2
XFILLER_168_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09332_ _09332_/A _09332_/B _09332_/C _10782_/A vssd1 vssd1 vccd1 vccd1 _09338_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_80_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_142_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09263_ _18980_/Q _18979_/Q _18978_/Q vssd1 vssd1 vccd1 vccd1 _09265_/C sky130_fd_sc_hd__or3_2
XFILLER_33_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_222_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09194_ _18569_/Q _18568_/Q _18567_/Q vssd1 vssd1 vccd1 vccd1 _09198_/A sky130_fd_sc_hd__or3_4
XFILLER_166_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_119_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_216_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_216_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_142_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08978_ _08979_/A vssd1 vssd1 vccd1 vccd1 _08978_/Y sky130_fd_sc_hd__inv_2
XFILLER_5_1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_229_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_216_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10940_ _10940_/A vssd1 vssd1 vccd1 vccd1 _10940_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_5_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_2_1_1_wb_clk_i clkbuf_2_1_1_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_3_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_205_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10871_ _10956_/A _10877_/B vssd1 vssd1 vccd1 vccd1 _10871_/X sky130_fd_sc_hd__or2_1
XFILLER_71_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_216_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_231_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12610_ _12618_/A _12610_/B vssd1 vssd1 vccd1 vccd1 _12612_/A sky130_fd_sc_hd__nor2_1
XPHY_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13590_ _18714_/Q _13581_/X _13582_/X _18708_/Q _13589_/X vssd1 vssd1 vccd1 vccd1
+ _13590_/X sky130_fd_sc_hd__a221o_1
XPHY_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_213_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12541_ _12574_/B _12542_/B vssd1 vssd1 vccd1 vccd1 _12556_/A sky130_fd_sc_hd__or2_1
XPHY_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_200_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15260_ _15301_/A _15263_/B vssd1 vssd1 vccd1 vccd1 _15260_/Y sky130_fd_sc_hd__nand2_1
XFILLER_196_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12472_ _12472_/A _12472_/B vssd1 vssd1 vccd1 vccd1 _12473_/A sky130_fd_sc_hd__and2_1
XFILLER_138_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_5_0_0_wb_clk_i clkbuf_5_1_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_5_0_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_2
X_14211_ _18209_/Q _14257_/B _14470_/A vssd1 vssd1 vccd1 vccd1 _14211_/X sky130_fd_sc_hd__o21a_1
XFILLER_138_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11423_ _11423_/A _12329_/B vssd1 vssd1 vccd1 vccd1 _11423_/Y sky130_fd_sc_hd__nand2_1
X_15191_ _15236_/A _15195_/B vssd1 vssd1 vccd1 vccd1 _15191_/Y sky130_fd_sc_hd__nand2_1
XFILLER_125_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14142_ _18371_/Q _13838_/X _14015_/A _18374_/Q _14141_/X vssd1 vssd1 vccd1 vccd1
+ _14142_/X sky130_fd_sc_hd__a221o_2
X_11354_ _13501_/A _11354_/B vssd1 vssd1 vccd1 vccd1 _11547_/B sky130_fd_sc_hd__xnor2_1
XFILLER_152_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10305_ _10301_/X _10304_/X _10305_/S vssd1 vssd1 vccd1 vccd1 _10312_/B sky130_fd_sc_hd__mux2_1
XFILLER_4_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_1319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14073_ _18842_/Q _13575_/X _13576_/X _18833_/Q _14072_/X vssd1 vssd1 vccd1 vccd1
+ _14073_/X sky130_fd_sc_hd__a221o_1
X_11285_ _11453_/A _11364_/A vssd1 vssd1 vccd1 vccd1 _11354_/B sky130_fd_sc_hd__nand2_1
X_18950_ _18950_/CLK _18950_/D vssd1 vssd1 vccd1 vccd1 _18950_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_140_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19059__30 vssd1 vssd1 vccd1 vccd1 _19059__30/HI _19153_/A sky130_fd_sc_hd__conb_1
X_10236_ _10236_/A vssd1 vssd1 vccd1 vccd1 _10236_/X sky130_fd_sc_hd__clkbuf_4
X_17901_ _17901_/CLK _17901_/D vssd1 vssd1 vccd1 vccd1 _17901_/Q sky130_fd_sc_hd__dfxtp_1
X_13024_ _17985_/Q _13015_/X _13023_/X vssd1 vssd1 vccd1 vccd1 _17985_/D sky130_fd_sc_hd__a21o_1
XFILLER_117_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18881_ _18914_/CLK _18881_/D vssd1 vssd1 vccd1 vccd1 _18881_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_121_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17832_ _18222_/CLK _17832_/D vssd1 vssd1 vccd1 vccd1 _17832_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_79_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10167_ _13009_/A _10167_/B vssd1 vssd1 vccd1 vccd1 _10170_/A sky130_fd_sc_hd__xor2_1
XFILLER_121_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17763_ _17763_/A vssd1 vssd1 vccd1 vccd1 _19024_/D sky130_fd_sc_hd__clkbuf_1
X_14975_ _14975_/A _15268_/B _14989_/C vssd1 vssd1 vccd1 vccd1 _14975_/X sky130_fd_sc_hd__or3_1
X_10098_ _09243_/A _10060_/X _10097_/X _09987_/A vssd1 vssd1 vccd1 vccd1 _10098_/X
+ sky130_fd_sc_hd__o211a_1
X_16714_ _16714_/A _16745_/B vssd1 vssd1 vccd1 vccd1 _16723_/B sky130_fd_sc_hd__nor2_2
XFILLER_212_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13926_ _18247_/Q _13715_/X _13513_/A _18241_/Q _13925_/X vssd1 vssd1 vccd1 vccd1
+ _13926_/X sky130_fd_sc_hd__a221o_1
XFILLER_48_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17694_ _17694_/A vssd1 vssd1 vccd1 vccd1 _18985_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_75_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_223_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16645_ _16648_/B _16642_/X _16644_/Y _16639_/X vssd1 vssd1 vccd1 vccd1 _18730_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_62_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13857_ _13857_/A vssd1 vssd1 vccd1 vccd1 _13858_/A sky130_fd_sc_hd__buf_8
XFILLER_35_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_228_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_1339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12808_ _12809_/A _17948_/Q vssd1 vssd1 vccd1 vccd1 _12808_/X sky130_fd_sc_hd__or2_1
X_16576_ _16575_/B _16574_/X _16575_/Y _16559_/X vssd1 vssd1 vccd1 vccd1 _18713_/D
+ sky130_fd_sc_hd__o211a_1
X_13788_ _18417_/Q _13651_/X _13783_/X _13787_/X vssd1 vssd1 vccd1 vccd1 _13788_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_37_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18315_ _18317_/CLK _18315_/D vssd1 vssd1 vccd1 vccd1 _18315_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_76_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15527_ _15527_/A _15599_/C vssd1 vssd1 vccd1 vccd1 _15534_/B sky130_fd_sc_hd__nor2_1
XFILLER_176_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_32_wb_clk_i clkbuf_5_7_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18809_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_12739_ _19002_/Q _19001_/Q _12739_/C _12948_/C vssd1 vssd1 vccd1 vccd1 _12742_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_176_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_188_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18246_ _18809_/CLK _18246_/D vssd1 vssd1 vccd1 vccd1 _18246_/Q sky130_fd_sc_hd__dfxtp_1
X_15458_ _18482_/Q _18446_/Q _15458_/S vssd1 vssd1 vccd1 vccd1 _15458_/X sky130_fd_sc_hd__mux2_1
XFILLER_175_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_204_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14409_ _18193_/Q _14409_/B vssd1 vssd1 vccd1 vccd1 _14414_/B sky130_fd_sc_hd__nor2_1
X_18177_ _18178_/CLK _18177_/D vssd1 vssd1 vccd1 vccd1 _18177_/Q sky130_fd_sc_hd__dfxtp_1
X_15389_ _15582_/A vssd1 vssd1 vccd1 vccd1 _15445_/A sky130_fd_sc_hd__clkbuf_2
X_17128_ _18844_/Q _17129_/B _17127_/Y _17117_/X vssd1 vssd1 vccd1 vccd1 _18844_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_183_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_1318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09950_ _10292_/S vssd1 vssd1 vccd1 vccd1 _09950_/X sky130_fd_sc_hd__buf_2
X_17059_ _17491_/A _17070_/B vssd1 vssd1 vccd1 vccd1 _17068_/B sky130_fd_sc_hd__nor2_1
XFILLER_100_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09881_ _09875_/A _09875_/B _09880_/X vssd1 vssd1 vccd1 vccd1 _09883_/B sky130_fd_sc_hd__a21bo_1
XFILLER_98_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_111_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_226_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_198_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_213_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09315_ _18464_/Q _18463_/Q _18462_/Q vssd1 vssd1 vccd1 vccd1 _09319_/A sky130_fd_sc_hd__or3_2
XFILLER_15_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_167_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09246_ _18896_/Q _18895_/Q _18894_/Q vssd1 vssd1 vccd1 vccd1 _09248_/C sky130_fd_sc_hd__or3_4
XFILLER_103_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09177_ _18593_/Q _18592_/Q _18591_/Q vssd1 vssd1 vccd1 vccd1 _09181_/A sky130_fd_sc_hd__or3_4
XFILLER_119_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_107_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_218_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11070_ _13442_/A vssd1 vssd1 vccd1 vccd1 _11070_/X sky130_fd_sc_hd__buf_2
XTAP_6025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10021_ _10940_/A _10017_/X _10020_/X _10010_/X vssd1 vssd1 vccd1 vccd1 _10021_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_6069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_193_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_229_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14760_ _14812_/A vssd1 vssd1 vccd1 vccd1 _14787_/S sky130_fd_sc_hd__clkbuf_2
XTAP_4689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11972_ _11932_/A _13438_/A _11946_/X _11948_/X vssd1 vssd1 vccd1 vccd1 _11973_/B
+ sky130_fd_sc_hd__a31o_1
XTAP_3955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13711_ _13699_/X _13709_/X _13710_/Y vssd1 vssd1 vccd1 vccd1 _13711_/X sky130_fd_sc_hd__o21a_2
XFILLER_205_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_189_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10923_ _10921_/X _10922_/X _10923_/S vssd1 vssd1 vccd1 vccd1 _10923_/X sky130_fd_sc_hd__mux2_1
XTAP_3988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14691_ _17747_/A vssd1 vssd1 vccd1 vccd1 _14778_/A sky130_fd_sc_hd__clkbuf_2
XTAP_3999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16430_ _16429_/B _16428_/X _16429_/Y _16418_/X vssd1 vssd1 vccd1 vccd1 _18677_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_186_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_189_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13642_ _13642_/A vssd1 vssd1 vccd1 vccd1 _13642_/X sky130_fd_sc_hd__buf_8
XFILLER_147_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10854_ _09360_/A _09365_/C _10870_/S vssd1 vssd1 vccd1 vccd1 _10854_/X sky130_fd_sc_hd__mux2_1
XFILLER_31_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16361_ _16389_/A _16364_/B vssd1 vssd1 vccd1 vccd1 _16361_/Y sky130_fd_sc_hd__nand2_1
XPHY_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_188_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13573_ _13573_/A vssd1 vssd1 vccd1 vccd1 _14081_/B sky130_fd_sc_hd__buf_6
XPHY_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10785_ _12099_/A _12100_/A vssd1 vssd1 vccd1 vccd1 _10843_/C sky130_fd_sc_hd__and2_2
XFILLER_125_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18100_ _18130_/CLK _18100_/D vssd1 vssd1 vccd1 vccd1 _18100_/Q sky130_fd_sc_hd__dfxtp_2
X_15312_ _15358_/A _15921_/B _15358_/C vssd1 vssd1 vccd1 vccd1 _15312_/X sky130_fd_sc_hd__or3_1
XFILLER_40_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_212_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12524_ _17916_/Q _17919_/Q vssd1 vssd1 vccd1 vccd1 _12535_/A sky130_fd_sc_hd__nand2b_2
XPHY_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16292_ _16325_/A _16294_/B vssd1 vssd1 vccd1 vccd1 _16292_/Y sky130_fd_sc_hd__nand2_1
XFILLER_188_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18031_ _18035_/CLK _18031_/D vssd1 vssd1 vccd1 vccd1 _18031_/Q sky130_fd_sc_hd__dfxtp_1
X_15243_ _15279_/A _15243_/B _15257_/C vssd1 vssd1 vccd1 vccd1 _15243_/X sky130_fd_sc_hd__or3_1
XFILLER_201_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12455_ _12455_/A vssd1 vssd1 vccd1 vccd1 _17903_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_185_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11406_ _11453_/A _11412_/A vssd1 vssd1 vccd1 vccd1 _11410_/A sky130_fd_sc_hd__xnor2_1
X_15174_ _15232_/A vssd1 vssd1 vccd1 vccd1 _15220_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_153_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12386_ _12388_/A _12388_/B _12388_/C vssd1 vssd1 vccd1 vccd1 _12397_/B sky130_fd_sc_hd__o21a_1
XFILLER_181_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14125_ _18899_/Q _14124_/X _13538_/A _18881_/Q vssd1 vssd1 vccd1 vccd1 _14125_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_207_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11337_ _11337_/A _12023_/B _11376_/A _11337_/D vssd1 vssd1 vccd1 vccd1 _11338_/A
+ sky130_fd_sc_hd__nand4_4
XFILLER_99_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_180_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_150_wb_clk_i clkbuf_5_27_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18373_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_141_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_125_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14056_ _18491_/Q _13619_/A _14052_/X _14055_/X vssd1 vssd1 vccd1 vccd1 _14056_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_45_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18933_ _18936_/CLK _18933_/D vssd1 vssd1 vccd1 vccd1 _18933_/Q sky130_fd_sc_hd__dfxtp_2
X_11268_ _13442_/A _13427_/A vssd1 vssd1 vccd1 vccd1 _11268_/Y sky130_fd_sc_hd__nor2_1
X_13007_ _13007_/A _13007_/B vssd1 vssd1 vccd1 vccd1 _13007_/Y sky130_fd_sc_hd__nand2_1
XFILLER_67_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10219_ _10215_/A _10215_/B _10218_/X vssd1 vssd1 vccd1 vccd1 _10220_/B sky130_fd_sc_hd__o21a_1
X_11199_ _11199_/A vssd1 vssd1 vccd1 vccd1 _17811_/D sky130_fd_sc_hd__clkbuf_1
X_18864_ _18866_/CLK _18864_/D vssd1 vssd1 vccd1 vccd1 _18864_/Q sky130_fd_sc_hd__dfxtp_2
X_17815_ _17821_/CLK _17815_/D vssd1 vssd1 vccd1 vccd1 _17815_/Q sky130_fd_sc_hd__dfxtp_1
X_18795_ _18812_/CLK _18795_/D vssd1 vssd1 vccd1 vccd1 _18795_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_5880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17746_ _17746_/A vssd1 vssd1 vccd1 vccd1 _19016_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_48_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14958_ _14958_/A vssd1 vssd1 vccd1 vccd1 _14974_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_130_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13909_ _18847_/Q _13735_/A _13734_/A _18853_/Q _13908_/X vssd1 vssd1 vccd1 vccd1
+ _13909_/X sky130_fd_sc_hd__a221o_1
XFILLER_47_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17677_ _14597_/A _17674_/Y _17675_/X _17676_/Y _18981_/Q vssd1 vssd1 vccd1 vccd1
+ _17678_/B sky130_fd_sc_hd__a32o_1
XINSDIODE2_210 _13562_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14889_ _14948_/A vssd1 vssd1 vccd1 vccd1 _14935_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_35_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XINSDIODE2_221 _13838_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XINSDIODE2_232 _17473_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16628_ _16678_/A _16773_/B _16628_/C vssd1 vssd1 vccd1 vccd1 _16628_/X sky130_fd_sc_hd__or3_1
XFILLER_23_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_243 _18316_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_189_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_254 _12027_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_265 _15175_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16559_ _16559_/A vssd1 vssd1 vccd1 vccd1 _16559_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_22_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_188_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09100_ _18794_/Q _18793_/Q _18792_/Q vssd1 vssd1 vccd1 vccd1 _09103_/B sky130_fd_sc_hd__or3_4
X_09031_ _09034_/A vssd1 vssd1 vccd1 vccd1 _09031_/Y sky130_fd_sc_hd__inv_2
XFILLER_176_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18229_ _18230_/CLK _18229_/D vssd1 vssd1 vccd1 vccd1 _18229_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_163_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_191_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_1262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_1295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09933_ _10348_/A vssd1 vssd1 vccd1 vccd1 _10292_/S sky130_fd_sc_hd__buf_2
XFILLER_131_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09864_ _18116_/Q _10113_/A vssd1 vssd1 vccd1 vccd1 _09867_/A sky130_fd_sc_hd__nand2_1
XFILLER_100_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09795_ _09812_/A _09812_/B vssd1 vssd1 vccd1 vccd1 _09795_/Y sky130_fd_sc_hd__nand2_1
XTAP_3207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_213_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_227_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_1277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_214_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_201_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_195_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10570_ _09294_/D _10568_/X _10569_/X _10036_/A vssd1 vssd1 vccd1 vccd1 _10570_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_50_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09229_ _18935_/Q _18934_/Q _18933_/Q vssd1 vssd1 vccd1 vccd1 _09232_/B sky130_fd_sc_hd__or3_2
XFILLER_166_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12240_ _12240_/A vssd1 vssd1 vccd1 vccd1 _17859_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_5_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_206_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12171_ _12170_/X _12171_/B _12171_/C vssd1 vssd1 vccd1 vccd1 _12171_/X sky130_fd_sc_hd__and3b_1
XFILLER_135_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_218_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11122_ _13452_/A _17808_/Q _11149_/S vssd1 vssd1 vccd1 vccd1 _11123_/A sky130_fd_sc_hd__mux2_1
XFILLER_174_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15930_ _15975_/A vssd1 vssd1 vccd1 vccd1 _15993_/B sky130_fd_sc_hd__buf_2
XFILLER_153_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11053_ _11895_/A vssd1 vssd1 vccd1 vccd1 _12272_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_49_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10004_ _10728_/A _10004_/B vssd1 vssd1 vccd1 vccd1 _10004_/X sky130_fd_sc_hd__or2_1
XFILLER_27_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15861_ _15925_/A vssd1 vssd1 vccd1 vccd1 _15861_/X sky130_fd_sc_hd__clkbuf_2
XTAP_4420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17600_ _17610_/A _17600_/B vssd1 vssd1 vccd1 vccd1 _17601_/A sky130_fd_sc_hd__and2_1
XTAP_5198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14812_ _14812_/A vssd1 vssd1 vccd1 vccd1 _14830_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_76_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18580_ _18593_/CLK _18580_/D vssd1 vssd1 vccd1 vccd1 _18580_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_4464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15792_ _15795_/B _15790_/X _15791_/Y _15783_/X vssd1 vssd1 vccd1 vccd1 _18526_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_188_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_224_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_229_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17531_ _17541_/A _17534_/B vssd1 vssd1 vccd1 vccd1 _17531_/Y sky130_fd_sc_hd__nand2_1
XTAP_3763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14743_ _14742_/B _14741_/X _14742_/Y _14738_/X vssd1 vssd1 vccd1 vccd1 _18275_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_29_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_229_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11955_ _11985_/A _11999_/B _11988_/A vssd1 vssd1 vccd1 vccd1 _11960_/C sky130_fd_sc_hd__and3_1
XTAP_3785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17462_ _17469_/B _17459_/X _17460_/X _17461_/X vssd1 vssd1 vccd1 vccd1 _18927_/D
+ sky130_fd_sc_hd__o211a_1
X_10906_ _14247_/A _12094_/A _10906_/C vssd1 vssd1 vccd1 vccd1 _10906_/X sky130_fd_sc_hd__or3_1
XFILLER_229_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14674_ _14687_/A _15266_/A vssd1 vssd1 vccd1 vccd1 _14683_/B sky130_fd_sc_hd__nor2_1
XFILLER_45_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11886_ _18160_/Q _11852_/X _11875_/Y vssd1 vssd1 vccd1 vccd1 _11887_/B sky130_fd_sc_hd__a21oi_1
XFILLER_220_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16413_ _18709_/Q _18673_/Q _16421_/S vssd1 vssd1 vccd1 vccd1 _16413_/X sky130_fd_sc_hd__mux2_1
X_19201_ _19201_/A _08985_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[1] sky130_fd_sc_hd__ebufn_8
X_13625_ _13841_/A vssd1 vssd1 vccd1 vccd1 _13625_/X sky130_fd_sc_hd__buf_8
X_17393_ _17395_/B _17391_/X _17392_/Y _17380_/X vssd1 vssd1 vccd1 vccd1 _18910_/D
+ sky130_fd_sc_hd__o211a_1
X_10837_ _09248_/A _09243_/A _09253_/B _10097_/A _10811_/A _10644_/A vssd1 vssd1 vccd1
+ vccd1 _10838_/C sky130_fd_sc_hd__mux4_1
XFILLER_160_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19132_ _19132_/A _09058_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[2] sky130_fd_sc_hd__ebufn_8
X_16344_ _16783_/A _16356_/B vssd1 vssd1 vccd1 vccd1 _16353_/B sky130_fd_sc_hd__nor2_2
XFILLER_186_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13556_ _18693_/Q _13551_/X _14014_/A _18696_/Q vssd1 vssd1 vccd1 vccd1 _13556_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_160_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10768_ _10768_/A vssd1 vssd1 vccd1 vccd1 _10768_/Y sky130_fd_sc_hd__inv_2
XFILLER_125_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_186_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12507_ _11767_/B _11761_/A _11767_/A vssd1 vssd1 vccd1 vccd1 _12528_/C sky130_fd_sc_hd__o21a_1
X_16275_ _16285_/B _16271_/X _16272_/X _16274_/X vssd1 vssd1 vccd1 vccd1 _18639_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_185_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13487_ _13563_/B _13541_/B vssd1 vssd1 vccd1 vccd1 _13652_/A sky130_fd_sc_hd__nor2_4
XFILLER_160_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10699_ _10818_/A vssd1 vssd1 vccd1 vccd1 _10700_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_218_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18014_ _18035_/CLK _18014_/D vssd1 vssd1 vccd1 vccd1 _18014_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_199_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15226_ _18431_/Q _18395_/Q _15226_/S vssd1 vssd1 vccd1 vccd1 _15226_/X sky130_fd_sc_hd__mux2_1
XFILLER_157_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12438_ _12419_/A _12439_/B _12439_/D _12439_/C vssd1 vssd1 vccd1 vccd1 _12438_/Y
+ sky130_fd_sc_hd__a31oi_2
XFILLER_201_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15157_ _16673_/A vssd1 vssd1 vccd1 vccd1 _15772_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_141_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12369_ _12472_/A _12369_/B _12369_/C vssd1 vssd1 vccd1 vccd1 _12370_/A sky130_fd_sc_hd__and3_1
XFILLER_141_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14108_ _18791_/Q _13524_/A _14106_/X _14107_/X vssd1 vssd1 vccd1 vccd1 _14108_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_153_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15088_ _15098_/A _15233_/B _15112_/C vssd1 vssd1 vccd1 vccd1 _15088_/X sky130_fd_sc_hd__or3_1
XFILLER_114_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14039_ _18323_/Q _13596_/A _13706_/X _18305_/Q vssd1 vssd1 vccd1 vccd1 _14039_/X
+ sky130_fd_sc_hd__a22o_1
X_18916_ _18931_/CLK _18916_/D vssd1 vssd1 vccd1 vccd1 _18916_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_113_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18847_ _18849_/CLK _18847_/D vssd1 vssd1 vccd1 vccd1 _18847_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_94_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_227_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09580_ _09580_/A _10705_/A vssd1 vssd1 vccd1 vccd1 _09580_/X sky130_fd_sc_hd__and2_1
XFILLER_67_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18778_ _18778_/CLK _18778_/D vssd1 vssd1 vccd1 vccd1 _18778_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_227_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17729_ _17729_/A vssd1 vssd1 vccd1 vccd1 _19008_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_70_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_208_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_189_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_1283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_1294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09014_ _09016_/A vssd1 vssd1 vccd1 vccd1 _09014_/Y sky130_fd_sc_hd__inv_2
XFILLER_192_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_117_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_219_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19113__84 vssd1 vssd1 vccd1 vccd1 _19113__84/HI _19221_/A sky130_fd_sc_hd__conb_1
XFILLER_137_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09916_ _09976_/A vssd1 vssd1 vccd1 vccd1 _09916_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_77_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_217_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09847_ _18126_/Q _09847_/B vssd1 vssd1 vccd1 vccd1 _09866_/A sky130_fd_sc_hd__xor2_4
XFILLER_100_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_1339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09778_ _09792_/A _09785_/B vssd1 vssd1 vccd1 vccd1 _09780_/B sky130_fd_sc_hd__xnor2_1
XTAP_3026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_215_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11740_ _11740_/A _11740_/B _11740_/C vssd1 vssd1 vccd1 vccd1 _11824_/A sky130_fd_sc_hd__nand3_2
XTAP_1624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_230_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11671_ _17861_/Q _11671_/B vssd1 vssd1 vccd1 vccd1 _11672_/B sky130_fd_sc_hd__nand2_1
XFILLER_35_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_1361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_169_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13410_ _13410_/A _13410_/B _13410_/C _13410_/D vssd1 vssd1 vccd1 vccd1 _13412_/A
+ sky130_fd_sc_hd__nor4_2
XFILLER_161_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10622_ _13007_/A _12102_/A vssd1 vssd1 vccd1 vccd1 _10622_/Y sky130_fd_sc_hd__nor2_1
X_14390_ _17640_/A vssd1 vssd1 vccd1 vccd1 _17564_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_127_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13341_ _18097_/Q _11042_/X _11025_/B _11045_/X _13339_/X vssd1 vssd1 vccd1 vccd1
+ _18097_/D sky130_fd_sc_hd__o221a_1
X_10553_ _10498_/A _10550_/X _10552_/X _10555_/A vssd1 vssd1 vccd1 vccd1 _10553_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_128_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_182_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16060_ _16115_/A _16666_/B _16115_/C vssd1 vssd1 vccd1 vccd1 _16060_/X sky130_fd_sc_hd__or3_1
XFILLER_194_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13272_ _13271_/Y _12951_/B _12927_/A _13269_/B vssd1 vssd1 vccd1 vccd1 _13272_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_108_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10484_ _10484_/A vssd1 vssd1 vccd1 vccd1 _10484_/X sky130_fd_sc_hd__buf_4
XFILLER_6_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_183_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15011_ _15252_/A vssd1 vssd1 vccd1 vccd1 _15061_/A sky130_fd_sc_hd__buf_2
XFILLER_6_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12223_ _17855_/Q _12222_/X _12233_/C vssd1 vssd1 vccd1 vccd1 _12223_/X sky130_fd_sc_hd__o21ba_1
XFILLER_123_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12154_ _13458_/A _12154_/B vssd1 vssd1 vccd1 vccd1 _12175_/B sky130_fd_sc_hd__or2_1
XFILLER_151_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11105_ _11719_/B vssd1 vssd1 vccd1 vccd1 _11720_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_151_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16962_ _16962_/A vssd1 vssd1 vccd1 vccd1 _17538_/B sky130_fd_sc_hd__buf_4
X_12085_ _12120_/A _12085_/B vssd1 vssd1 vccd1 vccd1 _12085_/Y sky130_fd_sc_hd__nor2_1
X_18701_ _18701_/CLK _18701_/D vssd1 vssd1 vccd1 vccd1 _18701_/Q sky130_fd_sc_hd__dfxtp_1
X_15913_ _15942_/A _15913_/B vssd1 vssd1 vccd1 vccd1 _15913_/Y sky130_fd_sc_hd__nand2_1
X_11036_ _11044_/A _11036_/B vssd1 vssd1 vccd1 vccd1 _13367_/A sky130_fd_sc_hd__nand2_1
X_16893_ _16999_/A vssd1 vssd1 vccd1 vccd1 _16893_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_209_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_231_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18632_ _18633_/CLK _18632_/D vssd1 vssd1 vccd1 vccd1 _18632_/Q sky130_fd_sc_hd__dfxtp_2
X_15844_ _15993_/A _15844_/B vssd1 vssd1 vccd1 vccd1 _15853_/B sky130_fd_sc_hd__nor2_1
XFILLER_37_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18563_ _18563_/CLK _18563_/D vssd1 vssd1 vccd1 vccd1 _18563_/Q sky130_fd_sc_hd__dfxtp_2
X_15775_ _18558_/Q _18522_/Q _15790_/S vssd1 vssd1 vccd1 vccd1 _15775_/X sky130_fd_sc_hd__mux2_1
XFILLER_224_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12987_ _12987_/A _13310_/A vssd1 vssd1 vccd1 vccd1 _12987_/Y sky130_fd_sc_hd__nand2_1
XTAP_3571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_220_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_206_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14726_ _14750_/A _14729_/B vssd1 vssd1 vccd1 vccd1 _14726_/Y sky130_fd_sc_hd__nand2_1
X_17514_ _17514_/A _17536_/B vssd1 vssd1 vccd1 vccd1 _17524_/B sky130_fd_sc_hd__nor2_2
X_18494_ _18496_/CLK _18494_/D vssd1 vssd1 vccd1 vccd1 _18494_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_205_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11938_ _11947_/A _11947_/B vssd1 vssd1 vccd1 vccd1 _12015_/A sky130_fd_sc_hd__nand2_2
XFILLER_60_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_1215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_220_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17445_ _17444_/B _17443_/X _17444_/Y _17441_/X vssd1 vssd1 vccd1 vccd1 _18923_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_2892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14657_ _18256_/Q _14658_/B _14656_/Y _14647_/X vssd1 vssd1 vccd1 vccd1 _18256_/D
+ sky130_fd_sc_hd__o211a_1
X_11869_ _11869_/A _11869_/B vssd1 vssd1 vccd1 vccd1 _11869_/Y sky130_fd_sc_hd__nand2_2
XFILLER_220_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13608_ _18840_/Q _13575_/A _13515_/X _18816_/Q _13607_/X vssd1 vssd1 vccd1 vccd1
+ _13608_/X sky130_fd_sc_hd__a221o_1
XFILLER_14_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17376_ _17376_/A _17516_/B _17376_/C vssd1 vssd1 vccd1 vccd1 _17376_/X sky130_fd_sc_hd__or3_1
XFILLER_158_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14588_ _18241_/Q _14589_/B _14586_/Y _14587_/X vssd1 vssd1 vccd1 vccd1 _18241_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_220_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16327_ _16327_/A vssd1 vssd1 vccd1 vccd1 _16345_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_203_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13539_ _13539_/A vssd1 vssd1 vccd1 vccd1 _13539_/X sky130_fd_sc_hd__buf_4
XFILLER_158_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_199_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16258_ _16701_/A _16307_/B vssd1 vssd1 vccd1 vccd1 _16268_/B sky130_fd_sc_hd__nor2_1
XFILLER_173_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_145_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15209_ _15206_/B _15205_/X _15206_/Y _15208_/X vssd1 vssd1 vccd1 vccd1 _18389_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_173_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16189_ _16188_/B _16187_/X _16188_/Y _16185_/X vssd1 vssd1 vccd1 vccd1 _18620_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_173_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_1366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_229_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_9 _09143_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09701_ _10036_/A vssd1 vssd1 vccd1 vccd1 _09987_/A sky130_fd_sc_hd__buf_2
XFILLER_101_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09632_ _17973_/Q vssd1 vssd1 vccd1 vccd1 _12946_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_228_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09563_ _09565_/A _09549_/B _09562_/X vssd1 vssd1 vccd1 vccd1 _09575_/A sky130_fd_sc_hd__a21oi_1
XFILLER_209_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09494_ _18191_/Q _18190_/Q _18189_/Q vssd1 vssd1 vccd1 vccd1 _09495_/B sky130_fd_sc_hd__or3_1
XFILLER_230_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_212_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_211_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_145_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_223_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_211_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_1348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_211_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_221_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_221_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_219_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_215_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_133_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_219_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12910_ _12913_/C _12910_/B vssd1 vssd1 vccd1 vccd1 _17966_/D sky130_fd_sc_hd__nor2_1
XFILLER_150_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13890_ _18985_/Q _14081_/B _13780_/X _18976_/Q _13889_/X vssd1 vssd1 vccd1 vccd1
+ _13890_/X sky130_fd_sc_hd__a221o_1
XFILLER_58_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12841_ _17945_/Q _17946_/Q vssd1 vssd1 vccd1 vccd1 _12843_/B sky130_fd_sc_hd__or2_1
XTAP_2100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_206_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15560_ _16005_/A _15597_/B vssd1 vssd1 vccd1 vccd1 _15570_/B sky130_fd_sc_hd__nor2_1
XTAP_1410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12772_ _13269_/B _12771_/Y _17941_/Q vssd1 vssd1 vccd1 vccd1 _12772_/Y sky130_fd_sc_hd__a21oi_1
XTAP_2155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_215_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14511_ _14511_/A vssd1 vssd1 vccd1 vccd1 _18227_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11723_ _17913_/Q vssd1 vssd1 vccd1 vccd1 _11753_/A sky130_fd_sc_hd__inv_2
XTAP_2199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15491_ _18489_/Q _18453_/Q _15494_/S vssd1 vssd1 vccd1 vccd1 _15491_/X sky130_fd_sc_hd__mux2_1
XTAP_1465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17230_ _17275_/A _17230_/B vssd1 vssd1 vccd1 vccd1 _17230_/Y sky130_fd_sc_hd__nand2_1
XFILLER_187_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14442_ _14422_/X _09503_/B _14423_/X vssd1 vssd1 vccd1 vccd1 _14442_/X sky130_fd_sc_hd__a21o_1
X_11654_ _11719_/B _11654_/B _11654_/C vssd1 vssd1 vccd1 vccd1 _11655_/C sky130_fd_sc_hd__and3_1
XFILLER_230_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10605_ _10605_/A _10605_/B _10605_/C _10605_/D vssd1 vssd1 vccd1 vccd1 _10897_/C
+ sky130_fd_sc_hd__and4_1
X_17161_ _17197_/A vssd1 vssd1 vccd1 vccd1 _17161_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_196_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14373_ _14373_/A _14373_/B _14373_/C vssd1 vssd1 vccd1 vccd1 _14373_/X sky130_fd_sc_hd__and3_1
X_11585_ _11661_/A _11499_/B _11261_/X _11501_/A _11584_/B vssd1 vssd1 vccd1 vccd1
+ _11587_/C sky130_fd_sc_hd__a2111oi_1
XFILLER_200_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_196_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16112_ _16714_/A _16150_/B vssd1 vssd1 vccd1 vccd1 _16123_/B sky130_fd_sc_hd__nor2_2
XFILLER_122_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13324_ _13324_/A _13324_/B vssd1 vssd1 vccd1 vccd1 _13324_/Y sky130_fd_sc_hd__nand2_1
XFILLER_196_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17092_ _17091_/B _17090_/X _17091_/Y _17076_/X vssd1 vssd1 vccd1 vccd1 _18836_/D
+ sky130_fd_sc_hd__o211a_1
X_10536_ _10935_/S _10536_/B vssd1 vssd1 vccd1 vccd1 _10536_/X sky130_fd_sc_hd__and2_1
XFILLER_6_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_155_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16043_ _16043_/A _16043_/B _16043_/C vssd1 vssd1 vccd1 vccd1 _16043_/X sky130_fd_sc_hd__or3_1
XFILLER_183_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13255_ _13255_/A _18082_/Q vssd1 vssd1 vccd1 vccd1 _13256_/A sky130_fd_sc_hd__and2_1
XFILLER_124_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10467_ _10463_/X _10465_/X _10902_/S vssd1 vssd1 vccd1 vccd1 _10467_/X sky130_fd_sc_hd__mux2_2
X_12206_ _11700_/Y _12205_/X _12205_/A _11704_/B vssd1 vssd1 vccd1 vccd1 _12207_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_108_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13186_ _13186_/A _18051_/Q vssd1 vssd1 vccd1 vccd1 _13187_/A sky130_fd_sc_hd__and2_1
X_10398_ _09916_/X _10396_/X _10397_/X _10278_/X vssd1 vssd1 vccd1 vccd1 _10399_/B
+ sky130_fd_sc_hd__a22oi_2
XFILLER_215_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12137_ _12151_/A vssd1 vssd1 vccd1 vccd1 _12158_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_17994_ _18108_/CLK _17994_/D vssd1 vssd1 vccd1 vccd1 _17994_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_96_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16945_ _16945_/A vssd1 vssd1 vccd1 vccd1 _17526_/A sky130_fd_sc_hd__buf_4
X_12068_ _12068_/A _13494_/B vssd1 vssd1 vccd1 vccd1 _12069_/D sky130_fd_sc_hd__xnor2_1
XFILLER_42_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11019_ _17972_/Q vssd1 vssd1 vccd1 vccd1 _11044_/A sky130_fd_sc_hd__inv_2
X_16876_ _17037_/A _16963_/C vssd1 vssd1 vccd1 vccd1 _16884_/B sky130_fd_sc_hd__nor2_2
XFILLER_133_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_231_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_226_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18615_ _18620_/CLK _18615_/D vssd1 vssd1 vccd1 vccd1 _18615_/Q sky130_fd_sc_hd__dfxtp_2
X_15827_ _18535_/Q _15829_/B _15826_/Y _15823_/X vssd1 vssd1 vccd1 vccd1 _18535_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_4080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_209_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15758_ _15821_/A vssd1 vssd1 vccd1 vccd1 _15894_/C sky130_fd_sc_hd__clkbuf_2
X_18546_ _18546_/CLK _18546_/D vssd1 vssd1 vccd1 vccd1 _18546_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_64_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_212_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_209_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14709_ _14772_/A vssd1 vssd1 vccd1 vccd1 _14841_/B sky130_fd_sc_hd__buf_2
X_15689_ _15694_/B _15686_/X _15688_/X _15681_/X vssd1 vssd1 vccd1 vccd1 _18501_/D
+ sky130_fd_sc_hd__o211a_1
X_18477_ _18482_/CLK _18477_/D vssd1 vssd1 vccd1 vccd1 _18477_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_53_1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17428_ _17453_/A _17432_/B vssd1 vssd1 vccd1 vccd1 _17428_/Y sky130_fd_sc_hd__nand2_1
XFILLER_220_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_1280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_220_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17359_ _18938_/Q _18902_/Q _17367_/S vssd1 vssd1 vccd1 vccd1 _17359_/X sky130_fd_sc_hd__mux2_1
XFILLER_88_1305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19029_ _19029_/CLK _19029_/D vssd1 vssd1 vccd1 vccd1 _19029_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_161_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_141_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08994_ _08997_/A vssd1 vssd1 vccd1 vccd1 _08994_/Y sky130_fd_sc_hd__inv_2
XFILLER_87_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_1330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_214_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_228_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_217_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09615_ _18117_/Q _18110_/Q vssd1 vssd1 vccd1 vccd1 _09617_/A sky130_fd_sc_hd__nand2_1
XFILLER_83_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09546_ _09544_/Y _09535_/B _09545_/Y vssd1 vssd1 vccd1 vccd1 _10142_/A sky130_fd_sc_hd__o21a_2
XFILLER_110_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09477_ _09474_/A _09463_/X _09461_/A _18142_/D vssd1 vssd1 vccd1 vccd1 _18141_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_212_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_141_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_180_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11370_ _11495_/B _11593_/B _11374_/C _11508_/C vssd1 vssd1 vccd1 vccd1 _11371_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_180_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10321_ _09277_/A _09277_/B _09277_/C _09277_/D _10307_/S _09905_/A vssd1 vssd1 vccd1
+ vccd1 _10321_/X sky130_fd_sc_hd__mux4_1
XFILLER_4_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13040_ _13009_/A _13025_/X _13039_/X _13037_/X vssd1 vssd1 vccd1 vccd1 _17992_/D
+ sky130_fd_sc_hd__o211a_1
X_10252_ _10206_/A _12074_/A _10251_/Y vssd1 vssd1 vccd1 vccd1 _11917_/A sky130_fd_sc_hd__a21o_1
XFILLER_191_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_1274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10183_ _10183_/A vssd1 vssd1 vccd1 vccd1 _10270_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_133_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14991_ _18373_/Q _18337_/Q _14994_/S vssd1 vssd1 vccd1 vccd1 _14991_/X sky130_fd_sc_hd__mux2_1
XFILLER_120_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16730_ _16752_/A _16732_/B vssd1 vssd1 vccd1 vccd1 _16730_/Y sky130_fd_sc_hd__nand2_1
X_13942_ _18784_/Q _13857_/A _13592_/A _18799_/Q _13941_/X vssd1 vssd1 vccd1 vccd1
+ _13942_/X sky130_fd_sc_hd__a221o_1
XFILLER_115_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16661_ _17265_/A _16976_/B vssd1 vssd1 vccd1 vccd1 _16727_/A sky130_fd_sc_hd__or2_1
XFILLER_74_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13873_ _18463_/Q _13581_/X _13871_/X _13872_/X vssd1 vssd1 vccd1 vccd1 _13873_/X
+ sky130_fd_sc_hd__a211o_1
Xclkbuf_leaf_175_wb_clk_i clkbuf_5_11_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18217_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_18400_ _18432_/CLK _18400_/D vssd1 vssd1 vccd1 vccd1 _18400_/Q sky130_fd_sc_hd__dfxtp_2
X_15612_ _15745_/B vssd1 vssd1 vccd1 vccd1 _15666_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_28_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12824_ _12824_/A vssd1 vssd1 vccd1 vccd1 _12824_/Y sky130_fd_sc_hd__inv_2
XFILLER_222_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16592_ _18753_/Q _18717_/Q _16598_/S vssd1 vssd1 vccd1 vccd1 _16592_/X sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_104_wb_clk_i clkbuf_5_28_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18582_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_222_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_216_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15543_ _15566_/A _15546_/B vssd1 vssd1 vccd1 vccd1 _15543_/Y sky130_fd_sc_hd__nand2_1
XFILLER_188_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18331_ _18343_/CLK _18331_/D vssd1 vssd1 vccd1 vccd1 _18331_/Q sky130_fd_sc_hd__dfxtp_2
X_12755_ _18017_/Q _18016_/Q _18019_/Q _18018_/Q vssd1 vssd1 vccd1 vccd1 _12920_/B
+ sky130_fd_sc_hd__and4_1
XTAP_1240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18262_ _18263_/CLK _18262_/D vssd1 vssd1 vccd1 vccd1 _18262_/Q sky130_fd_sc_hd__dfxtp_1
X_11706_ _11706_/A vssd1 vssd1 vccd1 vccd1 _11706_/Y sky130_fd_sc_hd__inv_2
XFILLER_15_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15474_ _15516_/A vssd1 vssd1 vccd1 vccd1 _15474_/X sky130_fd_sc_hd__buf_2
XFILLER_202_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12686_ _12685_/Y _17935_/Q _12697_/B _12676_/B vssd1 vssd1 vccd1 vccd1 _12686_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_147_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14425_ _18196_/Q _14424_/X _14401_/X _09499_/B vssd1 vssd1 vccd1 vccd1 _14426_/B
+ sky130_fd_sc_hd__o2bb2a_1
X_17213_ _17213_/A _17213_/B vssd1 vssd1 vccd1 vccd1 _17213_/Y sky130_fd_sc_hd__nand2_1
XFILLER_202_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11637_ _17861_/Q vssd1 vssd1 vccd1 vccd1 _11639_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_18193_ _18196_/CLK _18193_/D vssd1 vssd1 vccd1 vccd1 _18193_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_204_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_168_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_200_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17144_ _17143_/B _17142_/X _17143_/Y _17140_/X vssd1 vssd1 vccd1 vccd1 _18848_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_196_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14356_ _14354_/X _14272_/X _14355_/X _14340_/X vssd1 vssd1 vccd1 vccd1 _18182_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_204_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11568_ _11570_/A _12269_/A vssd1 vssd1 vccd1 vccd1 _11569_/B sky130_fd_sc_hd__nor2_1
XFILLER_183_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13307_ _18073_/Q _18072_/Q _18075_/Q _18074_/Q vssd1 vssd1 vccd1 vccd1 _13309_/B
+ sky130_fd_sc_hd__or4_1
XFILLER_6_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10519_ _09402_/B _09392_/D _09952_/A _09397_/A _10484_/A _10518_/X vssd1 vssd1 vccd1
+ vccd1 _10520_/B sky130_fd_sc_hd__mux4_2
X_17075_ _17088_/A _17080_/B vssd1 vssd1 vccd1 vccd1 _17075_/Y sky130_fd_sc_hd__nand2_1
XFILLER_115_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14287_ _14275_/X _14281_/X _14286_/X _14270_/X vssd1 vssd1 vccd1 vccd1 _18175_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_155_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11499_ _13509_/A _11499_/B _11499_/C _11922_/A vssd1 vssd1 vccd1 vccd1 _11499_/X
+ sky130_fd_sc_hd__and4b_1
XFILLER_226_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16026_ _18620_/Q _18584_/Q _16031_/S vssd1 vssd1 vccd1 vccd1 _16026_/X sky130_fd_sc_hd__mux2_1
XFILLER_143_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13238_ _13244_/A _18074_/Q vssd1 vssd1 vccd1 vccd1 _13239_/A sky130_fd_sc_hd__and2_1
XFILLER_100_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13169_ _13175_/A _18043_/Q vssd1 vssd1 vccd1 vccd1 _13170_/A sky130_fd_sc_hd__and2_1
XFILLER_151_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_170_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17977_ _19027_/CLK _17977_/D vssd1 vssd1 vccd1 vccd1 _17977_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_85_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16928_ _16928_/A vssd1 vssd1 vccd1 vccd1 _16947_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_111_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_225_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_226_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16859_ _18818_/Q _18782_/Q _16864_/S vssd1 vssd1 vccd1 vccd1 _16859_/X sky130_fd_sc_hd__mux2_1
XFILLER_65_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09400_ _18341_/Q _18340_/Q _18339_/Q vssd1 vssd1 vccd1 vccd1 _10877_/A sky130_fd_sc_hd__or3_2
XFILLER_0_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09331_ _18521_/Q _18520_/Q _18519_/Q vssd1 vssd1 vccd1 vccd1 _10782_/A sky130_fd_sc_hd__or3_4
X_18529_ _18533_/CLK _18529_/D vssd1 vssd1 vccd1 vccd1 _18529_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_34_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_222_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_221_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_209_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09262_ _18971_/Q _18970_/Q _18969_/Q vssd1 vssd1 vccd1 vccd1 _10813_/A sky130_fd_sc_hd__or3_2
XFILLER_205_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09193_ _09193_/A _09193_/B _09193_/C _09193_/D vssd1 vssd1 vccd1 vccd1 _09204_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_21_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_222_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_216_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_216_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08977_ _08979_/A vssd1 vssd1 vccd1 vccd1 _08977_/Y sky130_fd_sc_hd__inv_2
XTAP_4805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_2_wb_clk_i clkbuf_5_0_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17919_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_57_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_229_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_217_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_216_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_1207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10870_ _09413_/A _09418_/D _10870_/S vssd1 vssd1 vccd1 vccd1 _10870_/X sky130_fd_sc_hd__mux2_1
XFILLER_43_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_227_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_231_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09529_ _10113_/A _17784_/Q vssd1 vssd1 vccd1 vccd1 _09530_/B sky130_fd_sc_hd__or2_1
XFILLER_31_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12540_ _17921_/Q vssd1 vssd1 vccd1 vccd1 _12574_/B sky130_fd_sc_hd__inv_2
XPHY_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_196_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12471_ _12471_/A _12477_/D vssd1 vssd1 vccd1 vccd1 _12472_/B sky130_fd_sc_hd__xnor2_1
XFILLER_200_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_177_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14210_ _18208_/Q _14323_/C vssd1 vssd1 vccd1 vccd1 _14257_/B sky130_fd_sc_hd__and2_1
XFILLER_61_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11422_ _17881_/Q _17880_/Q vssd1 vssd1 vccd1 vccd1 _12329_/B sky130_fd_sc_hd__and2_1
X_15190_ _15247_/A vssd1 vssd1 vccd1 vccd1 _15236_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_165_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14141_ _18347_/Q _14017_/A _14137_/X _14140_/X vssd1 vssd1 vccd1 vccd1 _14141_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_125_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11353_ _11354_/B _11353_/B vssd1 vssd1 vccd1 vccd1 _11366_/A sky130_fd_sc_hd__and2_1
XFILLER_165_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10304_ _10278_/A _10302_/X _10303_/X _09976_/A vssd1 vssd1 vccd1 vccd1 _10304_/X
+ sky130_fd_sc_hd__a22o_1
X_14072_ _18815_/Q _13577_/X _14068_/X _14071_/X vssd1 vssd1 vccd1 vccd1 _14072_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_158_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11284_ _11359_/B _17799_/Q _17798_/Q vssd1 vssd1 vccd1 vccd1 _11364_/A sky130_fd_sc_hd__and3_2
XFILLER_98_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17900_ _17901_/CLK _17900_/D vssd1 vssd1 vccd1 vccd1 _17900_/Q sky130_fd_sc_hd__dfxtp_1
X_13023_ _13016_/X _12967_/A _12718_/X _11891_/X vssd1 vssd1 vccd1 vccd1 _13023_/X
+ sky130_fd_sc_hd__a31o_1
X_10235_ _10235_/A vssd1 vssd1 vccd1 vccd1 _10236_/A sky130_fd_sc_hd__buf_4
XFILLER_3_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18880_ _18914_/CLK _18880_/D vssd1 vssd1 vccd1 vccd1 _18880_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_121_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17831_ _18209_/CLK _17831_/D vssd1 vssd1 vccd1 vccd1 _17831_/Q sky130_fd_sc_hd__dfxtp_1
X_10166_ _10159_/A _10158_/A _10165_/X vssd1 vssd1 vccd1 vccd1 _10167_/B sky130_fd_sc_hd__a21bo_1
XFILLER_86_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19074__45 vssd1 vssd1 vccd1 vccd1 _19074__45/HI _19168_/A sky130_fd_sc_hd__conb_1
XFILLER_48_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17762_ _17764_/A _19025_/Q vssd1 vssd1 vccd1 vccd1 _17763_/A sky130_fd_sc_hd__and2_1
XFILLER_86_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14974_ _18369_/Q _18333_/Q _14974_/S vssd1 vssd1 vccd1 vccd1 _14974_/X sky130_fd_sc_hd__mux2_1
XFILLER_19_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10097_ _10097_/A _10103_/B vssd1 vssd1 vccd1 vccd1 _10097_/X sky130_fd_sc_hd__or2_1
XFILLER_43_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_208_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16713_ _16712_/B _16710_/X _16712_/Y _16704_/X vssd1 vssd1 vccd1 vccd1 _18746_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_207_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13925_ _18253_/Q _13716_/X _13490_/A _18244_/Q vssd1 vssd1 vccd1 vccd1 _13925_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_81_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17693_ _17712_/A _17693_/B vssd1 vssd1 vccd1 vccd1 _17694_/A sky130_fd_sc_hd__and2_1
XFILLER_208_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16644_ _16695_/A _16648_/B vssd1 vssd1 vccd1 vccd1 _16644_/Y sky130_fd_sc_hd__nand2_1
X_13856_ _13856_/A vssd1 vssd1 vccd1 vccd1 _13856_/X sky130_fd_sc_hd__buf_4
XFILLER_223_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12807_ _17921_/Q _17950_/Q vssd1 vssd1 vccd1 vccd1 _12807_/X sky130_fd_sc_hd__or2_1
XFILLER_34_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16575_ _16575_/A _16575_/B vssd1 vssd1 vccd1 vccd1 _16575_/Y sky130_fd_sc_hd__nand2_1
X_13787_ _18441_/Q _13663_/X _13784_/X _13786_/X vssd1 vssd1 vccd1 vccd1 _13787_/X
+ sky130_fd_sc_hd__a211o_1
X_10999_ _17821_/Q vssd1 vssd1 vccd1 vccd1 _11001_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_206_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18314_ _18317_/CLK _18314_/D vssd1 vssd1 vccd1 vccd1 _18314_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_37_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15526_ _15525_/B _15523_/X _15525_/Y _15516_/X vssd1 vssd1 vccd1 vccd1 _18461_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_204_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12738_ _18089_/Q _18000_/Q vssd1 vssd1 vccd1 vccd1 _12948_/C sky130_fd_sc_hd__and2b_2
XTAP_1081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15457_ _15460_/B _15454_/X _15456_/Y _15452_/X vssd1 vssd1 vccd1 vccd1 _18445_/D
+ sky130_fd_sc_hd__o211a_1
X_18245_ _18245_/CLK _18245_/D vssd1 vssd1 vccd1 vccd1 _18245_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_198_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12669_ _12665_/A _12665_/B _12663_/A vssd1 vssd1 vccd1 vccd1 _12672_/A sky130_fd_sc_hd__a21o_1
XFILLER_15_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14408_ _14420_/A _14408_/B vssd1 vssd1 vccd1 vccd1 _18192_/D sky130_fd_sc_hd__nor2_1
XFILLER_204_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15388_ _18467_/Q _18431_/Q _15388_/S vssd1 vssd1 vccd1 vccd1 _15388_/X sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_72_wb_clk_i clkbuf_5_23_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18650_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_198_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18176_ _18176_/CLK _18176_/D vssd1 vssd1 vccd1 vccd1 _18176_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_156_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17127_ _17152_/A _17129_/B vssd1 vssd1 vccd1 vccd1 _17127_/Y sky130_fd_sc_hd__nand2_1
X_14339_ _14299_/X _14282_/X _14283_/X _14300_/X _17119_/B vssd1 vssd1 vccd1 vccd1
+ _14339_/X sky130_fd_sc_hd__a311o_1
XFILLER_144_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17058_ _17056_/B _17055_/X _17056_/Y _17057_/X vssd1 vssd1 vccd1 vccd1 _18827_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_98_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16009_ _16017_/B _16006_/X _16007_/X _16008_/X vssd1 vssd1 vccd1 vccd1 _18579_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09880_ _09880_/A _09874_/A vssd1 vssd1 vccd1 vccd1 _09880_/X sky130_fd_sc_hd__or2b_1
XTAP_821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_214_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_213_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_202_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_210_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09314_ _09314_/A _09314_/B _09314_/C _09314_/D vssd1 vssd1 vccd1 vccd1 _09320_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_90_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_222_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_221_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09245_ _18908_/Q _18907_/Q _18906_/Q vssd1 vssd1 vccd1 vccd1 _09248_/B sky130_fd_sc_hd__or3_4
XFILLER_193_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_222_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09176_ _09176_/A _09176_/B _09176_/C _09176_/D vssd1 vssd1 vccd1 vccd1 _09187_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_147_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_116_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_6004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_116_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_6015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10020_ _10018_/X _10019_/X _10065_/A vssd1 vssd1 vccd1 vccd1 _10020_/X sky130_fd_sc_hd__mux2_1
XFILLER_49_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11971_ _12023_/B _11971_/B vssd1 vssd1 vccd1 vccd1 _13438_/A sky130_fd_sc_hd__nor2_2
XTAP_4679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13710_ _13710_/A _13710_/B _13710_/C vssd1 vssd1 vccd1 vccd1 _13710_/Y sky130_fd_sc_hd__nor3_4
XFILLER_229_1326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10922_ _09349_/A _09354_/A _09344_/A _09349_/B _10413_/A _10496_/A vssd1 vssd1 vccd1
+ vccd1 _10922_/X sky130_fd_sc_hd__mux4_1
XTAP_3978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14690_ _14734_/A _14690_/B _15279_/B vssd1 vssd1 vccd1 vccd1 _14690_/X sky130_fd_sc_hd__or3_1
XTAP_3989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13641_ _13735_/A vssd1 vssd1 vccd1 vccd1 _13642_/A sky130_fd_sc_hd__buf_8
XFILLER_32_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10853_ _09952_/A _09402_/B _09397_/A _09392_/D _14206_/A _10852_/X vssd1 vssd1 vccd1
+ vccd1 _10853_/X sky130_fd_sc_hd__mux4_1
XFILLER_112_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16360_ _18697_/Q _18661_/Q _16363_/S vssd1 vssd1 vccd1 vccd1 _16360_/X sky130_fd_sc_hd__mux2_1
XFILLER_125_1302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13572_ _13517_/X _13571_/X _12042_/B vssd1 vssd1 vccd1 vccd1 _13572_/X sky130_fd_sc_hd__o21a_2
XFILLER_38_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10784_ _10809_/A _10781_/X _10783_/X _10801_/S vssd1 vssd1 vccd1 vccd1 _10784_/X
+ sky130_fd_sc_hd__a211o_1
XPHY_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15311_ _16823_/A vssd1 vssd1 vccd1 vccd1 _15921_/B sky130_fd_sc_hd__buf_2
XFILLER_200_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_188_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12523_ _12635_/A vssd1 vssd1 vccd1 vccd1 _12523_/X sky130_fd_sc_hd__buf_2
XPHY_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16291_ _18642_/Q _16294_/B _16290_/X _16274_/X vssd1 vssd1 vccd1 vccd1 _18642_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_125_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_160_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_184_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_200_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15242_ _18435_/Q _18399_/Q _15246_/S vssd1 vssd1 vccd1 vccd1 _15242_/X sky130_fd_sc_hd__mux2_1
XFILLER_12_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18030_ _18030_/CLK _18030_/D vssd1 vssd1 vccd1 vccd1 _18030_/Q sky130_fd_sc_hd__dfxtp_1
X_19119__90 vssd1 vssd1 vccd1 vccd1 _19119__90/HI _19227_/A sky130_fd_sc_hd__conb_1
X_12454_ _12459_/A _12454_/B _12477_/A vssd1 vssd1 vccd1 vccd1 _12455_/A sky130_fd_sc_hd__and3_1
XFILLER_201_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11405_ _11405_/A _11656_/B vssd1 vssd1 vccd1 vccd1 _11732_/A sky130_fd_sc_hd__and2_2
X_15173_ _18417_/Q _18381_/Q _15177_/S vssd1 vssd1 vccd1 vccd1 _15173_/X sky130_fd_sc_hd__mux2_1
XFILLER_123_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12385_ _12397_/A _12385_/B vssd1 vssd1 vccd1 vccd1 _12388_/C sky130_fd_sc_hd__nor2_1
XFILLER_201_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14124_ _14124_/A vssd1 vssd1 vccd1 vccd1 _14124_/X sky130_fd_sc_hd__buf_8
XFILLER_153_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11336_ _11336_/A _11336_/B _11368_/B vssd1 vssd1 vccd1 vccd1 _11337_/D sky130_fd_sc_hd__or3b_1
XFILLER_181_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14055_ _18515_/Q _13837_/A _14053_/X _14054_/X vssd1 vssd1 vccd1 vccd1 _14055_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_84_1352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18932_ _18939_/CLK _18932_/D vssd1 vssd1 vccd1 vccd1 _18932_/Q sky130_fd_sc_hd__dfxtp_1
X_11267_ _11336_/B _11333_/A vssd1 vssd1 vccd1 vccd1 _11315_/B sky130_fd_sc_hd__nand2_1
XFILLER_97_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13006_ _12721_/X _13004_/X _13009_/B _12955_/X _17991_/Q vssd1 vssd1 vccd1 vccd1
+ _13006_/X sky130_fd_sc_hd__a32o_1
XFILLER_140_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10218_ _10218_/A _10218_/B vssd1 vssd1 vccd1 vccd1 _10218_/X sky130_fd_sc_hd__or2_1
X_18863_ _18865_/CLK _18863_/D vssd1 vssd1 vccd1 vccd1 _18863_/Q sky130_fd_sc_hd__dfxtp_4
X_11198_ _11205_/C _11198_/B _11198_/C vssd1 vssd1 vccd1 vccd1 _11199_/A sky130_fd_sc_hd__and3b_1
XFILLER_132_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_190_wb_clk_i clkbuf_5_9_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18157_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_45_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_1339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17814_ _18989_/CLK _17814_/D vssd1 vssd1 vccd1 vccd1 _17814_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_94_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10149_ _10175_/A _10175_/B _10147_/A _10178_/A vssd1 vssd1 vccd1 vccd1 _10172_/A
+ sky130_fd_sc_hd__a211o_1
XFILLER_212_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18794_ _18812_/CLK _18794_/D vssd1 vssd1 vccd1 vccd1 _18794_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_43_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17745_ _17745_/A _19017_/Q vssd1 vssd1 vccd1 vccd1 _17746_/A sky130_fd_sc_hd__and2_1
XFILLER_54_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14957_ _14960_/B _14955_/X _14956_/Y _14941_/X vssd1 vssd1 vccd1 vccd1 _18328_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_82_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13908_ _18856_/Q _13489_/A _13763_/A _18871_/Q vssd1 vssd1 vccd1 vccd1 _13908_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_36_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_200 _11820_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17676_ _17674_/Y _17631_/A _14386_/A vssd1 vssd1 vccd1 vccd1 _17676_/Y sky130_fd_sc_hd__a21oi_1
X_14888_ _18347_/Q _18311_/Q _14905_/S vssd1 vssd1 vccd1 vccd1 _14888_/X sky130_fd_sc_hd__mux2_1
XINSDIODE2_211 _13580_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_222 _14064_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16627_ _16808_/A vssd1 vssd1 vccd1 vccd1 _16678_/A sky130_fd_sc_hd__dlymetal6s2s_1
XINSDIODE2_233 _14977_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13839_ _18694_/Q _13838_/X _13612_/A _18697_/Q vssd1 vssd1 vccd1 vccd1 _13839_/X
+ sky130_fd_sc_hd__a22o_1
XINSDIODE2_244 _18326_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_255 _13492_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XINSDIODE2_266 _17265_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16558_ _16572_/A _16562_/B vssd1 vssd1 vccd1 vccd1 _16558_/Y sky130_fd_sc_hd__nand2_1
XFILLER_91_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15509_ _15511_/B _15507_/X _15508_/Y _15496_/X vssd1 vssd1 vccd1 vccd1 _18457_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_175_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16489_ _16783_/A _16501_/B vssd1 vssd1 vccd1 vccd1 _16499_/B sky130_fd_sc_hd__nor2_2
XFILLER_176_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09030_ _09034_/A vssd1 vssd1 vccd1 vccd1 _09030_/Y sky130_fd_sc_hd__inv_2
XFILLER_176_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18228_ _18230_/CLK _18228_/D vssd1 vssd1 vccd1 vccd1 _18228_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_191_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_191_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18159_ _18209_/CLK _18159_/D vssd1 vssd1 vccd1 vccd1 _18159_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_89_1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_1274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_137_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09932_ _09932_/A _09932_/B vssd1 vssd1 vccd1 vccd1 _09932_/X sky130_fd_sc_hd__or2_1
XFILLER_132_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_207_wb_clk_i clkbuf_5_6_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18970_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09863_ _18116_/Q _18112_/Q vssd1 vssd1 vccd1 vccd1 _09867_/B sky130_fd_sc_hd__or2_1
XFILLER_86_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09794_ _09787_/A _09787_/B _09793_/X vssd1 vssd1 vccd1 vccd1 _09812_/B sky130_fd_sc_hd__o21a_1
XFILLER_6_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_227_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_1272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_213_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_214_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_210_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09228_ _18950_/Q _18949_/Q _18948_/Q vssd1 vssd1 vccd1 vccd1 _10826_/A sky130_fd_sc_hd__or3_4
XFILLER_194_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_182_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09159_ _18662_/Q _18661_/Q _18660_/Q vssd1 vssd1 vccd1 vccd1 _09160_/D sky130_fd_sc_hd__or3_4
XFILLER_182_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12170_ _12158_/A _12168_/X _12180_/A vssd1 vssd1 vccd1 vccd1 _12170_/X sky130_fd_sc_hd__o21ba_1
XFILLER_107_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_194_1366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11121_ _11895_/A vssd1 vssd1 vccd1 vccd1 _11149_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_150_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11052_ _12217_/A vssd1 vssd1 vccd1 vccd1 _11895_/A sky130_fd_sc_hd__buf_2
XFILLER_231_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10003_ _09114_/A _09119_/B _10003_/S vssd1 vssd1 vccd1 vccd1 _10003_/X sky130_fd_sc_hd__mux2_1
XFILLER_131_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15860_ _15873_/A _15865_/B vssd1 vssd1 vccd1 vccd1 _15860_/Y sky130_fd_sc_hd__nand2_1
XTAP_4410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19044__15 vssd1 vssd1 vccd1 vccd1 _19044__15/HI _19138_/A sky130_fd_sc_hd__conb_1
XTAP_4432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14811_ _14814_/B _14809_/X _14810_/Y _14799_/X vssd1 vssd1 vccd1 vccd1 _18292_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_97_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15791_ _15815_/A _15795_/B vssd1 vssd1 vccd1 vccd1 _15791_/Y sky130_fd_sc_hd__nand2_1
XTAP_4465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_218_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17530_ _18982_/Q _18946_/Q _17533_/S vssd1 vssd1 vccd1 vccd1 _17530_/X sky130_fd_sc_hd__mux2_1
XTAP_4498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14742_ _14753_/A _14742_/B vssd1 vssd1 vccd1 vccd1 _14742_/Y sky130_fd_sc_hd__nand2_1
X_11954_ _12041_/B _11961_/B vssd1 vssd1 vccd1 vccd1 _11988_/A sky130_fd_sc_hd__or2_2
XTAP_3764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10905_ _09386_/A _09376_/B _09381_/C _09972_/A _12089_/A _10852_/X vssd1 vssd1 vccd1
+ vccd1 _10906_/C sky130_fd_sc_hd__mux4_1
XFILLER_189_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14673_ _16945_/A vssd1 vssd1 vccd1 vccd1 _15266_/A sky130_fd_sc_hd__buf_6
XFILLER_60_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17461_ _17497_/A vssd1 vssd1 vccd1 vccd1 _17461_/X sky130_fd_sc_hd__clkbuf_2
X_11885_ _12207_/A _11885_/B vssd1 vssd1 vccd1 vccd1 _17834_/D sky130_fd_sc_hd__nor2_1
XFILLER_225_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_229_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19200_ _19200_/A _09059_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[0] sky130_fd_sc_hd__ebufn_8
X_16412_ _16417_/B _16410_/X _16411_/X _16398_/X vssd1 vssd1 vccd1 vccd1 _18672_/D
+ sky130_fd_sc_hd__o211a_1
X_13624_ _13624_/A vssd1 vssd1 vccd1 vccd1 _13841_/A sky130_fd_sc_hd__buf_6
XFILLER_177_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10836_ _10689_/A _10835_/X _10766_/A vssd1 vssd1 vccd1 vccd1 _10836_/X sky130_fd_sc_hd__a21o_1
X_17392_ _17392_/A _17395_/B vssd1 vssd1 vccd1 vccd1 _17392_/Y sky130_fd_sc_hd__nand2_1
XFILLER_73_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19131_ _19131_/A _09057_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[1] sky130_fd_sc_hd__ebufn_8
XFILLER_201_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16343_ _16342_/B _16340_/X _16342_/Y _16334_/X vssd1 vssd1 vccd1 vccd1 _18656_/D
+ sky130_fd_sc_hd__o211a_1
X_13555_ _13573_/A vssd1 vssd1 vccd1 vccd1 _14014_/A sky130_fd_sc_hd__buf_2
XFILLER_13_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_186_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10767_ _09176_/A _09176_/C _09186_/D _09181_/B _10662_/A _10812_/S vssd1 vssd1 vccd1
+ vccd1 _10768_/A sky130_fd_sc_hd__mux4_2
XFILLER_34_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_125_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_158_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12506_ _17519_/A vssd1 vssd1 vccd1 vccd1 _17427_/S sky130_fd_sc_hd__buf_2
X_16274_ _16354_/A vssd1 vssd1 vccd1 vccd1 _16274_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_173_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13486_ _17803_/Q _13509_/B vssd1 vssd1 vccd1 vccd1 _13541_/B sky130_fd_sc_hd__nand2b_4
X_10698_ _10801_/S vssd1 vssd1 vccd1 vccd1 _10818_/A sky130_fd_sc_hd__buf_2
XFILLER_200_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15225_ _15227_/B _15222_/X _15223_/Y _15224_/X vssd1 vssd1 vccd1 vccd1 _18394_/D
+ sky130_fd_sc_hd__o211a_1
X_18013_ _18035_/CLK _18013_/D vssd1 vssd1 vccd1 vccd1 _18013_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_218_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12437_ _12437_/A _12437_/B vssd1 vssd1 vccd1 vccd1 _12439_/C sky130_fd_sc_hd__or2_1
XFILLER_154_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_201_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15156_ _15156_/A _15279_/C vssd1 vssd1 vccd1 vccd1 _15169_/B sky130_fd_sc_hd__nor2_1
XFILLER_160_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12368_ _12365_/X _12366_/X _12353_/A vssd1 vssd1 vccd1 vccd1 _12369_/C sky130_fd_sc_hd__a21o_1
XFILLER_99_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14107_ _18797_/Q _13697_/A _13598_/X _18773_/Q vssd1 vssd1 vccd1 vccd1 _14107_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_126_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11319_ _17877_/Q vssd1 vssd1 vccd1 vccd1 _11323_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_15087_ _18396_/Q _18360_/Q _15100_/S vssd1 vssd1 vccd1 vccd1 _15087_/X sky130_fd_sc_hd__mux2_1
XFILLER_4_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12299_ _17879_/Q _12299_/B _12299_/C vssd1 vssd1 vccd1 vccd1 _12300_/B sky130_fd_sc_hd__or3_1
XFILLER_45_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14038_ _18326_/Q _13561_/A _13492_/A _18317_/Q vssd1 vssd1 vccd1 vccd1 _14038_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_80_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18915_ _18931_/CLK _18915_/D vssd1 vssd1 vccd1 vccd1 _18915_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_86_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18846_ _18871_/CLK _18846_/D vssd1 vssd1 vccd1 vccd1 _18846_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_110_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_227_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18777_ _18778_/CLK _18777_/D vssd1 vssd1 vccd1 vccd1 _18777_/Q sky130_fd_sc_hd__dfxtp_2
X_15989_ _15991_/B _15986_/X _15987_/Y _15988_/X vssd1 vssd1 vccd1 vccd1 _18574_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_224_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17728_ _17734_/A _19009_/Q vssd1 vssd1 vccd1 vccd1 _17729_/A sky130_fd_sc_hd__and2_1
XFILLER_24_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_224_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17659_ _17659_/A _17659_/B vssd1 vssd1 vccd1 vccd1 _17660_/A sky130_fd_sc_hd__and2_1
XFILLER_211_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_177_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09013_ _09016_/A vssd1 vssd1 vccd1 vccd1 _09013_/Y sky130_fd_sc_hd__inv_2
XFILLER_128_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_176_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_219_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09915_ _09915_/A _12130_/A vssd1 vssd1 vccd1 vccd1 _09976_/A sky130_fd_sc_hd__nor2_2
XFILLER_28_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_217_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_219_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09846_ _09846_/A _09846_/B vssd1 vssd1 vccd1 vccd1 _09847_/B sky130_fd_sc_hd__nand2_1
XTAP_470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_224_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09777_ _09777_/A vssd1 vssd1 vccd1 vccd1 _10213_/A sky130_fd_sc_hd__buf_2
XTAP_3016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_226_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11670_ _11648_/X _11653_/B _11848_/B _11666_/Y _11669_/X vssd1 vssd1 vccd1 vccd1
+ _11670_/X sky130_fd_sc_hd__o41a_1
XFILLER_199_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_148_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_230_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10621_ _10705_/A _10706_/B vssd1 vssd1 vccd1 vccd1 _12102_/A sky130_fd_sc_hd__xor2_4
XFILLER_139_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_224_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_195_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13340_ _18096_/Q _13336_/X _13337_/X _13339_/X vssd1 vssd1 vccd1 vccd1 _18096_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_210_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10552_ _10561_/S _10552_/B vssd1 vssd1 vccd1 vccd1 _10552_/X sky130_fd_sc_hd__and2b_1
XFILLER_168_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13271_ _13271_/A vssd1 vssd1 vccd1 vccd1 _13271_/Y sky130_fd_sc_hd__inv_2
XFILLER_182_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10483_ _09114_/B _09109_/B _09119_/C _09109_/C _10413_/A _10454_/X vssd1 vssd1 vccd1
+ vccd1 _10483_/X sky130_fd_sc_hd__mux4_2
Xclkbuf_leaf_129_wb_clk_i clkbuf_5_24_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18392_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_33_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15010_ _15649_/A vssd1 vssd1 vccd1 vccd1 _15252_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_185_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12222_ _17858_/Q _11602_/B _17859_/Q vssd1 vssd1 vccd1 vccd1 _12222_/X sky130_fd_sc_hd__a21o_1
XFILLER_142_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_151_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12153_ _17841_/Q _12171_/B _12152_/X _11863_/X vssd1 vssd1 vccd1 vccd1 _17841_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_151_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11104_ _11466_/B vssd1 vssd1 vccd1 vccd1 _11719_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_190_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16961_ _18840_/Q _18804_/Q _16970_/S vssd1 vssd1 vccd1 vccd1 _16961_/X sky130_fd_sc_hd__mux2_1
X_12084_ _12084_/A _12084_/B vssd1 vssd1 vccd1 vccd1 _12085_/B sky130_fd_sc_hd__xnor2_4
XFILLER_1_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18700_ _18701_/CLK _18700_/D vssd1 vssd1 vccd1 vccd1 _18700_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_150_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15912_ _18556_/Q _15913_/B _15911_/Y _15901_/X vssd1 vssd1 vccd1 vccd1 _18556_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_42_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11035_ _13368_/B _11035_/B vssd1 vssd1 vccd1 vccd1 _13398_/A sky130_fd_sc_hd__or2_1
X_16892_ _17323_/A vssd1 vssd1 vccd1 vccd1 _16999_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_65_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18631_ _18633_/CLK _18631_/D vssd1 vssd1 vccd1 vccd1 _18631_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_209_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15843_ _15839_/B _15838_/X _15839_/Y _15842_/X vssd1 vssd1 vccd1 vccd1 _18539_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_4240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18562_ _18572_/CLK _18562_/D vssd1 vssd1 vccd1 vccd1 _18562_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_218_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15774_ _15863_/A vssd1 vssd1 vccd1 vccd1 _15790_/S sky130_fd_sc_hd__clkbuf_2
XTAP_4295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12986_ _13000_/C vssd1 vssd1 vccd1 vccd1 _12990_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_206_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17513_ _17512_/B _17511_/X _17512_/Y _17497_/X vssd1 vssd1 vccd1 vccd1 _18941_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_91_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14725_ _18307_/Q _18271_/Q _14736_/S vssd1 vssd1 vccd1 vccd1 _14725_/X sky130_fd_sc_hd__mux2_1
XFILLER_79_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18493_ _18497_/CLK _18493_/D vssd1 vssd1 vccd1 vccd1 _18493_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_3594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11937_ _11934_/Y _11944_/A _11937_/C _11984_/B vssd1 vssd1 vccd1 vccd1 _11937_/X
+ sky130_fd_sc_hd__and4bb_1
XFILLER_73_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17444_ _17456_/A _17444_/B vssd1 vssd1 vccd1 vccd1 _17444_/Y sky130_fd_sc_hd__nand2_1
XTAP_2893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14656_ _14681_/A _14658_/B vssd1 vssd1 vccd1 vccd1 _14656_/Y sky130_fd_sc_hd__nand2_1
X_11868_ _11869_/A _11868_/B vssd1 vssd1 vccd1 vccd1 _11868_/X sky130_fd_sc_hd__or2_1
XFILLER_177_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_1298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13607_ _18822_/Q _13568_/X _13605_/X _13606_/X vssd1 vssd1 vccd1 vccd1 _13607_/X
+ sky130_fd_sc_hd__a211o_1
X_10819_ _10833_/A _10819_/B _10910_/D _10819_/D vssd1 vssd1 vccd1 vccd1 _10822_/C
+ sky130_fd_sc_hd__and4_1
XFILLER_220_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17375_ _18942_/Q _18906_/Q _17386_/S vssd1 vssd1 vccd1 vccd1 _17375_/X sky130_fd_sc_hd__mux2_1
XFILLER_186_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14587_ _14668_/A vssd1 vssd1 vccd1 vccd1 _14587_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_14_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11799_ _11781_/Y _11783_/Y _11784_/X _11763_/X _11798_/X vssd1 vssd1 vccd1 vccd1
+ _11799_/X sky130_fd_sc_hd__a221o_1
XFILLER_229_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16326_ _16329_/B _16324_/X _16325_/Y _16314_/X vssd1 vssd1 vccd1 vccd1 _18652_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_9_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_199_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13538_ _13538_/A vssd1 vssd1 vccd1 vccd1 _13539_/A sky130_fd_sc_hd__buf_6
XFILLER_173_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_203_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_199_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16257_ _16256_/B _16255_/X _16256_/Y _16252_/X vssd1 vssd1 vccd1 vccd1 _18635_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_146_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13469_ _14421_/A vssd1 vssd1 vccd1 vccd1 _13480_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_64_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15208_ _15283_/A vssd1 vssd1 vccd1 vccd1 _15208_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_145_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16188_ _16202_/A _16188_/B vssd1 vssd1 vccd1 vccd1 _16188_/Y sky130_fd_sc_hd__nand2_1
XFILLER_142_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15139_ _15178_/A _15142_/B vssd1 vssd1 vccd1 vccd1 _15139_/Y sky130_fd_sc_hd__nand2_1
XFILLER_47_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_114_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09700_ _10024_/A vssd1 vssd1 vccd1 vccd1 _10036_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_68_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09631_ _09645_/A _09631_/B vssd1 vssd1 vccd1 vccd1 _09637_/A sky130_fd_sc_hd__xnor2_1
X_18829_ _18858_/CLK _18829_/D vssd1 vssd1 vccd1 vccd1 _18829_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_67_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_1322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09562_ _09580_/A _10618_/A vssd1 vssd1 vccd1 vccd1 _09562_/X sky130_fd_sc_hd__and2_1
XFILLER_167_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_1340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_224_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09493_ _14383_/A vssd1 vssd1 vccd1 vccd1 _17591_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_212_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_168_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_212_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_1232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_222_wb_clk_i _17803_/CLK vssd1 vssd1 vccd1 vccd1 _17806_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_219_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_180_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_219_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_191_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_219_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_219_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09829_ _11032_/A _09834_/B _09828_/X vssd1 vssd1 vccd1 vccd1 _12112_/B sky130_fd_sc_hd__a21o_1
XFILLER_100_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12840_ _12840_/A vssd1 vssd1 vccd1 vccd1 _17945_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_74_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_230_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_215_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12771_ _13318_/A _12769_/Y _12770_/Y vssd1 vssd1 vccd1 vccd1 _12771_/Y sky130_fd_sc_hd__o21ai_1
XTAP_1400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_215_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_199_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11722_ _11727_/A vssd1 vssd1 vccd1 vccd1 _11767_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_14510_ _17556_/A _14510_/B _14510_/C vssd1 vssd1 vccd1 vccd1 _14511_/A sky130_fd_sc_hd__and3_1
XTAP_2178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15490_ _15931_/A _15548_/B vssd1 vssd1 vccd1 vccd1 _15500_/B sky130_fd_sc_hd__nor2_1
XFILLER_203_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11653_ _11653_/A _11653_/B vssd1 vssd1 vccd1 vccd1 _11653_/Y sky130_fd_sc_hd__nand2_1
XFILLER_35_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14441_ _14441_/A vssd1 vssd1 vccd1 vccd1 _18200_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_120_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_161_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_230_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10604_ _12126_/A _10598_/X _10602_/X _09889_/A _10603_/X vssd1 vssd1 vccd1 vccd1
+ _10605_/D sky130_fd_sc_hd__a32o_1
XFILLER_11_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14372_ _14507_/A _14372_/B vssd1 vssd1 vccd1 vccd1 _14373_/B sky130_fd_sc_hd__nor2_1
X_17160_ _17193_/A _17449_/B _17173_/C vssd1 vssd1 vccd1 vccd1 _17160_/X sky130_fd_sc_hd__or3_1
XFILLER_31_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11584_ _11784_/A _11584_/B _11784_/B vssd1 vssd1 vccd1 vccd1 _11783_/A sky130_fd_sc_hd__and3_1
XFILLER_196_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16111_ _16862_/A vssd1 vssd1 vccd1 vccd1 _16714_/A sky130_fd_sc_hd__buf_8
XFILLER_122_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13323_ _13329_/B _13322_/Y _13318_/X vssd1 vssd1 vccd1 vccd1 _13324_/B sky130_fd_sc_hd__a21o_1
XFILLER_6_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_196_1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10535_ _09695_/X _09696_/X _09697_/X _09698_/X _10561_/S _10503_/S vssd1 vssd1 vccd1
+ vccd1 _10536_/B sky130_fd_sc_hd__mux4_2
XFILLER_122_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17091_ _17091_/A _17091_/B vssd1 vssd1 vccd1 vccd1 _17091_/Y sky130_fd_sc_hd__nand2_1
XFILLER_13_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16042_ _18624_/Q _18588_/Q _16050_/S vssd1 vssd1 vccd1 vccd1 _16042_/X sky130_fd_sc_hd__mux2_1
XFILLER_129_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13254_ _13254_/A vssd1 vssd1 vccd1 vccd1 _18080_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_109_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10466_ _10466_/A vssd1 vssd1 vccd1 vccd1 _10902_/S sky130_fd_sc_hd__buf_4
XFILLER_136_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12205_ _12205_/A _12210_/B vssd1 vssd1 vccd1 vccd1 _12205_/X sky130_fd_sc_hd__and2_1
X_13185_ _13185_/A vssd1 vssd1 vccd1 vccd1 _18049_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_123_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10397_ _09248_/B _09243_/B _09253_/C _09243_/C _09971_/S _09923_/X vssd1 vssd1 vccd1
+ vccd1 _10397_/X sky130_fd_sc_hd__mux4_1
Xclkbuf_3_6_0_wb_clk_i clkbuf_3_7_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_6_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_151_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12136_ _17944_/Q _18168_/Q _12144_/S vssd1 vssd1 vccd1 vccd1 _12151_/A sky130_fd_sc_hd__mux2_2
XFILLER_97_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17993_ _18061_/CLK _17993_/D vssd1 vssd1 vccd1 vccd1 _17993_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_215_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16944_ _16943_/B _16942_/X _16943_/Y _16940_/X vssd1 vssd1 vccd1 vccd1 _18800_/D
+ sky130_fd_sc_hd__o211a_1
X_12067_ _12067_/A _12067_/B _12066_/Y vssd1 vssd1 vccd1 vccd1 _12069_/C sky130_fd_sc_hd__or3b_1
Xclkbuf_leaf_97_wb_clk_i clkbuf_5_18_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18263_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_38_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11018_ _11018_/A vssd1 vssd1 vccd1 vccd1 _11018_/Y sky130_fd_sc_hd__inv_2
XFILLER_42_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16875_ _16874_/B _16873_/X _16874_/Y _16871_/X vssd1 vssd1 vccd1 vccd1 _18785_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_42_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_26_wb_clk_i clkbuf_5_6_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18936_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_37_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_225_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_231_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18614_ _18614_/CLK _18614_/D vssd1 vssd1 vccd1 vccd1 _18614_/Q sky130_fd_sc_hd__dfxtp_2
X_15826_ _15873_/A _15829_/B vssd1 vssd1 vccd1 vccd1 _15826_/Y sky130_fd_sc_hd__nand2_1
XTAP_4070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_225_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18545_ _18557_/CLK _18545_/D vssd1 vssd1 vccd1 vccd1 _18545_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_92_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15757_ _15757_/A _17549_/A vssd1 vssd1 vccd1 vccd1 _15821_/A sky130_fd_sc_hd__or2_1
XTAP_3380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12969_ _12969_/A _12969_/B _12969_/C vssd1 vssd1 vccd1 vccd1 _12970_/B sky130_fd_sc_hd__nor3_1
XFILLER_221_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14708_ _15292_/A _14843_/C vssd1 vssd1 vccd1 vccd1 _14715_/B sky130_fd_sc_hd__nor2_2
XFILLER_209_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18476_ _18482_/CLK _18476_/D vssd1 vssd1 vccd1 vccd1 _18476_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_221_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15688_ _15734_/A _15984_/B _15724_/C vssd1 vssd1 vccd1 vccd1 _15688_/X sky130_fd_sc_hd__or3_1
XFILLER_21_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_220_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17427_ _18955_/Q _18919_/Q _17427_/S vssd1 vssd1 vccd1 vccd1 _17427_/X sky130_fd_sc_hd__mux2_1
X_14639_ _14651_/A _15229_/A vssd1 vssd1 vccd1 vccd1 _14646_/B sky130_fd_sc_hd__nor2_1
XFILLER_18_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_221_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_221_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_1292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_220_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17358_ _17360_/B _17356_/X _17357_/Y _17341_/X vssd1 vssd1 vccd1 vccd1 _18901_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_158_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16309_ _18684_/Q _18648_/Q _16324_/S vssd1 vssd1 vccd1 vccd1 _16309_/X sky130_fd_sc_hd__mux2_1
XFILLER_118_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17289_ _18920_/Q _18884_/Q _17298_/S vssd1 vssd1 vccd1 vccd1 _17289_/X sky130_fd_sc_hd__mux2_1
XFILLER_101_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19028_ _19028_/CLK _19028_/D vssd1 vssd1 vccd1 vccd1 _19028_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_173_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_216_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08993_ _08997_/A vssd1 vssd1 vccd1 vccd1 _08993_/Y sky130_fd_sc_hd__inv_2
XFILLER_138_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_228_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_1304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_228_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_217_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09614_ _18117_/Q _18110_/Q vssd1 vssd1 vccd1 vccd1 _09617_/B sky130_fd_sc_hd__or2_1
XFILLER_44_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09545_ _18097_/Q _13000_/C vssd1 vssd1 vccd1 vccd1 _09545_/Y sky130_fd_sc_hd__nand2_1
XFILLER_225_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_224_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_1271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09476_ _09474_/Y _09482_/B _18138_/D vssd1 vssd1 vccd1 vccd1 _18140_/D sky130_fd_sc_hd__o21a_1
XFILLER_180_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_197_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_212_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10320_ _14260_/B _10315_/X _10319_/X _10605_/B vssd1 vssd1 vccd1 vccd1 _10320_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_109_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10251_ _10253_/A _10829_/A _13348_/A vssd1 vssd1 vccd1 vccd1 _10251_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_191_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10182_ _10456_/A _10438_/A vssd1 vssd1 vccd1 vccd1 _10183_/A sky130_fd_sc_hd__and2_4
XFILLER_191_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14990_ _14995_/B _14986_/X _14989_/X _14980_/X vssd1 vssd1 vccd1 vccd1 _18336_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_8_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13941_ _18793_/Q _13716_/X _13579_/A _18787_/Q vssd1 vssd1 vccd1 vccd1 _13941_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_120_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16660_ _16658_/B _16657_/X _16658_/Y _16659_/X vssd1 vssd1 vccd1 vccd1 _18734_/D
+ sky130_fd_sc_hd__o211a_1
X_13872_ _18472_/Q _13531_/A _13598_/X _18448_/Q vssd1 vssd1 vccd1 vccd1 _13872_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_75_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_207_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15611_ _15677_/A vssd1 vssd1 vccd1 vccd1 _15745_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_216_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12823_ _12530_/Y _17945_/Q _12815_/Y _12662_/B _12822_/X vssd1 vssd1 vccd1 vccd1
+ _12823_/X sky130_fd_sc_hd__a221o_1
X_16591_ _16734_/A _16602_/B vssd1 vssd1 vccd1 vccd1 _16599_/B sky130_fd_sc_hd__nor2_1
XFILLER_34_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18330_ _18346_/CLK _18330_/D vssd1 vssd1 vccd1 vccd1 _18330_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_43_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15542_ _18502_/Q _18466_/Q _15545_/S vssd1 vssd1 vccd1 vccd1 _15542_/X sky130_fd_sc_hd__mux2_1
XFILLER_188_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12754_ _18011_/Q _18010_/Q _12948_/C _12754_/D vssd1 vssd1 vccd1 vccd1 _12920_/A
+ sky130_fd_sc_hd__and4_1
XTAP_1241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_231_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18261_ _18263_/CLK _18261_/D vssd1 vssd1 vccd1 vccd1 _18261_/Q sky130_fd_sc_hd__dfxtp_1
X_11705_ _11698_/X _11702_/X _11705_/C _11705_/D vssd1 vssd1 vccd1 vccd1 _11705_/X
+ sky130_fd_sc_hd__and4bb_1
XTAP_1274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15473_ _15511_/A _15473_/B vssd1 vssd1 vccd1 vccd1 _15473_/Y sky130_fd_sc_hd__nand2_1
XTAP_1285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12685_ _12697_/B _12676_/B _17932_/Q vssd1 vssd1 vccd1 vccd1 _12685_/Y sky130_fd_sc_hd__o21ai_1
XTAP_1296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_144_wb_clk_i clkbuf_5_26_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18278_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_42_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17212_ _18902_/Q _18866_/Q _17221_/S vssd1 vssd1 vccd1 vccd1 _17212_/X sky130_fd_sc_hd__mux2_1
XFILLER_24_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11636_ _11620_/Y _11631_/X _11635_/X vssd1 vssd1 vccd1 vccd1 _11680_/C sky130_fd_sc_hd__a21oi_1
X_14424_ _14422_/X _09498_/B _14423_/X vssd1 vssd1 vccd1 vccd1 _14424_/X sky130_fd_sc_hd__a21o_1
XFILLER_198_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18192_ _18991_/CLK _18192_/D vssd1 vssd1 vccd1 vccd1 _18192_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_11_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17143_ _17156_/A _17143_/B vssd1 vssd1 vccd1 vccd1 _17143_/Y sky130_fd_sc_hd__nand2_1
X_11567_ _17866_/Q _17865_/Q vssd1 vssd1 vccd1 vccd1 _11570_/A sky130_fd_sc_hd__nor2_1
X_14355_ _17942_/Q _14355_/B _14355_/C _14355_/D vssd1 vssd1 vccd1 vccd1 _14355_/X
+ sky130_fd_sc_hd__or4_1
XFILLER_200_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10518_ _10518_/A vssd1 vssd1 vccd1 vccd1 _10518_/X sky130_fd_sc_hd__buf_2
X_13306_ _18077_/Q _18076_/Q _18079_/Q _18078_/Q vssd1 vssd1 vccd1 vccd1 _13309_/A
+ sky130_fd_sc_hd__or4_1
XFILLER_143_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17074_ _18868_/Q _18832_/Q _17074_/S vssd1 vssd1 vccd1 vccd1 _17074_/X sky130_fd_sc_hd__mux2_1
X_14286_ _14243_/X _14282_/X _14283_/X _14244_/X _15145_/B vssd1 vssd1 vccd1 vccd1
+ _14286_/X sky130_fd_sc_hd__a311o_1
XFILLER_144_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11498_ _11498_/A _11541_/A vssd1 vssd1 vccd1 vccd1 _11499_/C sky130_fd_sc_hd__and2_1
X_16025_ _16027_/B _16023_/X _16024_/Y _16008_/X vssd1 vssd1 vccd1 vccd1 _18583_/D
+ sky130_fd_sc_hd__o211a_1
X_13237_ _13237_/A vssd1 vssd1 vccd1 vccd1 _18072_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_226_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10449_ _10550_/S vssd1 vssd1 vccd1 vccd1 _10450_/S sky130_fd_sc_hd__buf_4
XFILLER_97_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13168_ _13168_/A vssd1 vssd1 vccd1 vccd1 _18041_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_152_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_123_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12119_ _12119_/A _12119_/B vssd1 vssd1 vccd1 vccd1 _14267_/B sky130_fd_sc_hd__xnor2_4
XFILLER_111_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13099_ _13107_/A _18011_/Q vssd1 vssd1 vccd1 vccd1 _13100_/A sky130_fd_sc_hd__and2_1
X_17976_ _18108_/CLK _17976_/D vssd1 vssd1 vccd1 vccd1 _17976_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_69_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16927_ _16930_/B _16925_/X _16926_/Y _16917_/X vssd1 vssd1 vccd1 vccd1 _18796_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_37_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16858_ _16860_/B _16856_/X _16857_/Y _16848_/X vssd1 vssd1 vccd1 vccd1 _18781_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_93_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_226_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15809_ _18567_/Q _18531_/Q _15809_/S vssd1 vssd1 vccd1 vccd1 _15809_/X sky130_fd_sc_hd__mux2_1
XFILLER_81_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_1310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_207_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16789_ _16813_/A _16792_/B vssd1 vssd1 vccd1 vccd1 _16789_/Y sky130_fd_sc_hd__nand2_1
XFILLER_225_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_209_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_209_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09330_ _18536_/Q _18535_/Q _18534_/Q vssd1 vssd1 vccd1 vccd1 _09332_/C sky130_fd_sc_hd__or3_4
X_18528_ _18533_/CLK _18528_/D vssd1 vssd1 vccd1 vccd1 _18528_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_20_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09261_ _18977_/Q _18976_/Q _18975_/Q vssd1 vssd1 vccd1 vccd1 _09265_/A sky130_fd_sc_hd__or3_2
XFILLER_222_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18459_ _18467_/CLK _18459_/D vssd1 vssd1 vccd1 vccd1 _18459_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_181_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09192_ _18590_/Q _18589_/Q _18588_/Q vssd1 vssd1 vccd1 vccd1 _09193_/D sky130_fd_sc_hd__or3_2
XFILLER_222_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08976_ _08979_/A vssd1 vssd1 vccd1 vccd1 _08976_/Y sky130_fd_sc_hd__inv_2
XFILLER_88_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_217_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_229_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_217_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_205_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09528_ _10113_/A _17784_/Q vssd1 vssd1 vccd1 vccd1 _09530_/A sky130_fd_sc_hd__nand2_1
XPHY_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_231_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_213_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09459_ _09467_/A vssd1 vssd1 vccd1 vccd1 _18138_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_24_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_227_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_212_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_184_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12470_ _17906_/Q _12470_/B vssd1 vssd1 vccd1 vccd1 _12477_/D sky130_fd_sc_hd__xor2_1
XFILLER_71_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_131_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_229_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11421_ _17881_/Q _17880_/Q vssd1 vssd1 vccd1 vccd1 _12323_/A sky130_fd_sc_hd__or2_1
XFILLER_137_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14140_ _18359_/Q _14124_/X _14138_/X _14139_/X vssd1 vssd1 vccd1 vccd1 _14140_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_137_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11352_ _11392_/B _11364_/A vssd1 vssd1 vccd1 vccd1 _11353_/B sky130_fd_sc_hd__or2_1
XFILLER_4_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10303_ _09219_/A _09209_/C _10795_/A _09214_/C _10376_/B _09937_/A vssd1 vssd1 vccd1
+ vccd1 _10303_/X sky130_fd_sc_hd__mux4_1
XFILLER_4_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14071_ _18839_/Q _13551_/X _14069_/X _14070_/X vssd1 vssd1 vccd1 vccd1 _14071_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_180_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11283_ _11869_/A vssd1 vssd1 vccd1 vccd1 _11820_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_193_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13022_ _12958_/A _13015_/X _13021_/X _13011_/X vssd1 vssd1 vccd1 vccd1 _17984_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_112_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_180_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10234_ _10542_/A vssd1 vssd1 vccd1 vccd1 _10235_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_152_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17830_ _18217_/CLK _17830_/D vssd1 vssd1 vccd1 vccd1 _17830_/Q sky130_fd_sc_hd__dfxtp_1
X_10165_ _10158_/A _10159_/A _10165_/S vssd1 vssd1 vccd1 vccd1 _10165_/X sky130_fd_sc_hd__mux2_1
XFILLER_121_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17761_ _17761_/A vssd1 vssd1 vccd1 vccd1 _19023_/D sky130_fd_sc_hd__clkbuf_1
X_14973_ _15266_/A _14985_/B vssd1 vssd1 vccd1 vccd1 _14983_/B sky130_fd_sc_hd__nor2_2
X_10096_ _09248_/A _09253_/B _10096_/S vssd1 vssd1 vccd1 vccd1 _10096_/X sky130_fd_sc_hd__mux2_1
XFILLER_47_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_208_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16712_ _16755_/A _16712_/B vssd1 vssd1 vccd1 vccd1 _16712_/Y sky130_fd_sc_hd__nand2_1
X_13924_ _13637_/Y _13883_/X _13915_/X _13923_/X vssd1 vssd1 vccd1 vccd1 _13924_/X
+ sky130_fd_sc_hd__a211o_2
XFILLER_208_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17692_ _17641_/X _17687_/Y _17675_/X _17688_/Y _18985_/Q vssd1 vssd1 vccd1 vccd1
+ _17693_/B sky130_fd_sc_hd__a32o_1
XFILLER_75_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16643_ _16828_/A vssd1 vssd1 vccd1 vccd1 _16695_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_78_1349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13855_ _18733_/Q _13575_/X _13576_/X _18724_/Q _13854_/X vssd1 vssd1 vccd1 vccd1
+ _13855_/X sky130_fd_sc_hd__a221o_2
XFILLER_207_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12806_ _17921_/Q _17950_/Q vssd1 vssd1 vccd1 vccd1 _12806_/Y sky130_fd_sc_hd__nand2_1
XFILLER_90_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16574_ _18749_/Q _18713_/Q _16598_/S vssd1 vssd1 vccd1 vccd1 _16574_/X sky130_fd_sc_hd__mux2_1
XFILLER_204_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13786_ _18429_/Q _13785_/X _13766_/X _18411_/Q vssd1 vssd1 vccd1 vccd1 _13786_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_16_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10998_ _17820_/Q vssd1 vssd1 vccd1 vccd1 _11232_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_204_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18313_ _18317_/CLK _18313_/D vssd1 vssd1 vccd1 vccd1 _18313_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_31_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15525_ _15570_/A _15525_/B vssd1 vssd1 vccd1 vccd1 _15525_/Y sky130_fd_sc_hd__nand2_1
XFILLER_204_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_5_27_0_wb_clk_i clkbuf_5_27_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_5_27_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_2
XTAP_1071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12737_ _19004_/Q _19003_/Q _19006_/Q _19005_/Q vssd1 vssd1 vccd1 vccd1 _12739_/C
+ sky130_fd_sc_hd__and4_1
XFILLER_31_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_203_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18244_ _18244_/CLK _18244_/D vssd1 vssd1 vccd1 vccd1 _18244_/Q sky130_fd_sc_hd__dfxtp_1
X_15456_ _15508_/A _15460_/B vssd1 vssd1 vccd1 vccd1 _15456_/Y sky130_fd_sc_hd__nand2_1
XFILLER_176_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12668_ _12662_/B _12635_/X _12665_/Y _12666_/X _12667_/X vssd1 vssd1 vccd1 vccd1
+ _17931_/D sky130_fd_sc_hd__a221o_1
XFILLER_30_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14407_ _18192_/Q _14406_/X _14401_/X _14409_/B vssd1 vssd1 vccd1 vccd1 _14408_/B
+ sky130_fd_sc_hd__o2bb2a_1
X_11619_ _11619_/A vssd1 vssd1 vccd1 vccd1 _11619_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_30_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18175_ _18178_/CLK _18175_/D vssd1 vssd1 vccd1 vccd1 _18175_/Q sky130_fd_sc_hd__dfxtp_1
X_15387_ _15390_/B _15384_/X _15386_/Y _15382_/X vssd1 vssd1 vccd1 vccd1 _18430_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_204_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_190_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12599_ _17926_/Q _12594_/B _12582_/A _12582_/B _12589_/A vssd1 vssd1 vccd1 vccd1
+ _12600_/C sky130_fd_sc_hd__o221ai_4
XFILLER_128_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17126_ _18843_/Q _17129_/B _17125_/X _17117_/X vssd1 vssd1 vccd1 vccd1 _18843_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_156_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14338_ _18179_/Q vssd1 vssd1 vccd1 vccd1 _17119_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_183_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17057_ _17096_/A vssd1 vssd1 vccd1 vccd1 _17057_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_144_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14269_ _14243_/X _14227_/X _14229_/X _14244_/X _18173_/Q vssd1 vssd1 vccd1 vccd1
+ _14269_/X sky130_fd_sc_hd__a311o_1
XFILLER_83_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16008_ _16028_/A vssd1 vssd1 vccd1 vccd1 _16008_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_83_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_41_wb_clk_i _18759_/CLK vssd1 vssd1 vccd1 vccd1 _18764_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_124_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17959_ _17959_/CLK _17959_/D vssd1 vssd1 vccd1 vccd1 _17959_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_22_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_226_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_122_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_214_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_213_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_213_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09313_ _18473_/Q _18472_/Q _18471_/Q vssd1 vssd1 vccd1 vccd1 _09314_/D sky130_fd_sc_hd__or3_4
XFILLER_22_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_210_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_222_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09244_ _18893_/Q _18892_/Q _18891_/Q vssd1 vssd1 vccd1 vccd1 _09248_/A sky130_fd_sc_hd__or3_4
XFILLER_221_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09175_ _18596_/Q _18595_/Q _18594_/Q vssd1 vssd1 vccd1 vccd1 _09176_/D sky130_fd_sc_hd__or3_2
XFILLER_119_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_222_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_6005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_227_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_1272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08959_ _08960_/A vssd1 vssd1 vccd1 vccd1 _08959_/Y sky130_fd_sc_hd__inv_2
XTAP_4625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_229_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11970_ _11970_/A _11975_/A _11970_/C vssd1 vssd1 vccd1 vccd1 _11971_/B sky130_fd_sc_hd__nor3_1
XTAP_3935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10921_ _09344_/B _09354_/C _10391_/A _10389_/A _10484_/X _10231_/X vssd1 vssd1 vccd1
+ vccd1 _10921_/X sky130_fd_sc_hd__mux4_1
XTAP_3968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_229_1338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13640_ _13677_/A vssd1 vssd1 vccd1 vccd1 _13735_/A sky130_fd_sc_hd__buf_6
XFILLER_16_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10852_ _10852_/A vssd1 vssd1 vccd1 vccd1 _10852_/X sky130_fd_sc_hd__buf_4
XFILLER_32_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_201_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13571_ _18681_/Q _13525_/X _13540_/X _13570_/X vssd1 vssd1 vccd1 vccd1 _13571_/X
+ sky130_fd_sc_hd__a211o_1
X_10783_ _09327_/A _10781_/S _10782_/X _10668_/A vssd1 vssd1 vccd1 vccd1 _10783_/X
+ sky130_fd_sc_hd__o211a_1
XPHY_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_227_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15310_ _18450_/Q _18414_/Q _15334_/S vssd1 vssd1 vccd1 vccd1 _15310_/X sky130_fd_sc_hd__mux2_1
XFILLER_213_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_1268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_201_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_197_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12522_ _12522_/A vssd1 vssd1 vccd1 vccd1 _12635_/A sky130_fd_sc_hd__clkbuf_2
XPHY_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16290_ _16310_/A _16880_/B _16333_/C vssd1 vssd1 vccd1 vccd1 _16290_/X sky130_fd_sc_hd__or3_1
XFILLER_188_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_201_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15241_ _15241_/A _15277_/B vssd1 vssd1 vccd1 vccd1 _15253_/B sky130_fd_sc_hd__nor2_2
XFILLER_200_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12453_ _12452_/A _12452_/B _12452_/C vssd1 vssd1 vccd1 vccd1 _12477_/A sky130_fd_sc_hd__a21o_1
XFILLER_172_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11404_ _11404_/A _11404_/B vssd1 vssd1 vccd1 vccd1 _11656_/B sky130_fd_sc_hd__nand2_1
XFILLER_201_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15172_ _15172_/A _15229_/B vssd1 vssd1 vccd1 vccd1 _15182_/B sky130_fd_sc_hd__nor2_2
XFILLER_153_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12384_ _17895_/Q _12384_/B _12384_/C vssd1 vssd1 vccd1 vccd1 _12385_/B sky130_fd_sc_hd__nor3_1
XFILLER_197_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11335_ _11333_/Y _11334_/X _11301_/A vssd1 vssd1 vccd1 vccd1 _11376_/A sky130_fd_sc_hd__a21oi_4
X_14123_ _18884_/Q _14019_/X _13500_/X _18908_/Q vssd1 vssd1 vccd1 vccd1 _14123_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_21_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18931_ _18931_/CLK _18931_/D vssd1 vssd1 vccd1 vccd1 _18931_/Q sky130_fd_sc_hd__dfxtp_1
X_14054_ _18503_/Q _14124_/A _13706_/X _18485_/Q vssd1 vssd1 vccd1 vccd1 _14054_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_10_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11266_ _11764_/A _11770_/B _11254_/Y _11265_/X vssd1 vssd1 vccd1 vccd1 _11905_/A
+ sky130_fd_sc_hd__a31o_2
XFILLER_113_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13005_ _13005_/A _13005_/B vssd1 vssd1 vccd1 vccd1 _13009_/B sky130_fd_sc_hd__nand2_1
X_10217_ _10217_/A _10217_/B vssd1 vssd1 vccd1 vccd1 _10221_/B sky130_fd_sc_hd__xnor2_2
XFILLER_140_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18862_ _18862_/CLK _18862_/D vssd1 vssd1 vccd1 vccd1 _18862_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_171_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11197_ _11196_/B _11190_/A _11196_/D _17811_/Q vssd1 vssd1 vccd1 vccd1 _11198_/C
+ sky130_fd_sc_hd__a31o_1
XFILLER_67_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17813_ _18989_/CLK _17813_/D vssd1 vssd1 vccd1 vccd1 _17813_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_121_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10148_ _10144_/A _10148_/B vssd1 vssd1 vccd1 vccd1 _10178_/A sky130_fd_sc_hd__and2b_1
X_18793_ _18823_/CLK _18793_/D vssd1 vssd1 vccd1 vccd1 _18793_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17744_ _17744_/A vssd1 vssd1 vccd1 vccd1 _19015_/D sky130_fd_sc_hd__clkbuf_1
XTAP_5893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14956_ _14992_/A _14960_/B vssd1 vssd1 vccd1 vccd1 _14956_/Y sky130_fd_sc_hd__nand2_1
X_10079_ _09227_/C _09232_/B _09237_/D _09232_/D _10955_/S _10065_/A vssd1 vssd1 vccd1
+ vccd1 _10079_/X sky130_fd_sc_hd__mux4_1
XFILLER_63_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_169_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13907_ _18874_/Q _13657_/X _13544_/A _18850_/Q _13906_/X vssd1 vssd1 vccd1 vccd1
+ _13907_/X sky130_fd_sc_hd__a221o_1
XFILLER_223_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17675_ _17675_/A vssd1 vssd1 vccd1 vccd1 _17675_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_169_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14887_ _14958_/A vssd1 vssd1 vccd1 vccd1 _14905_/S sky130_fd_sc_hd__clkbuf_2
XINSDIODE2_201 _12207_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XINSDIODE2_212 _13585_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16626_ _18762_/Q _18726_/Q _16637_/S vssd1 vssd1 vccd1 vccd1 _16626_/X sky130_fd_sc_hd__mux2_1
XINSDIODE2_223 _14436_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13838_ _13838_/A vssd1 vssd1 vccd1 vccd1 _13838_/X sky130_fd_sc_hd__buf_6
XFILLER_35_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_234 _17228_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_245 _17449_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_256 _13575_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_267 _16666_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16557_ _18745_/Q _18709_/Q _16565_/S vssd1 vssd1 vccd1 vccd1 _16557_/X sky130_fd_sc_hd__mux2_1
XFILLER_50_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13769_ _18489_/Q _13733_/X _13762_/X _13768_/X vssd1 vssd1 vccd1 vccd1 _13769_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_50_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15508_ _15508_/A _15511_/B vssd1 vssd1 vccd1 vccd1 _15508_/Y sky130_fd_sc_hd__nand2_1
X_16488_ _16487_/B _16486_/X _16487_/Y _16477_/X vssd1 vssd1 vccd1 vccd1 _18692_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_31_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18227_ _18230_/CLK _18227_/D vssd1 vssd1 vccd1 vccd1 _18227_/Q sky130_fd_sc_hd__dfxtp_1
X_15439_ _15445_/B _15435_/X _15438_/X _15428_/X vssd1 vssd1 vccd1 vccd1 _18441_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_15_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_106_1280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18158_ _18163_/CLK _18158_/D vssd1 vssd1 vccd1 vccd1 hold4/A sky130_fd_sc_hd__dfxtp_1
XFILLER_8_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17109_ _17136_/A _17538_/B _17109_/C vssd1 vssd1 vccd1 vccd1 _17109_/X sky130_fd_sc_hd__or3_1
XFILLER_116_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18089_ _18993_/CLK _18089_/D vssd1 vssd1 vccd1 vccd1 _18089_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_102_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09931_ _09921_/X _09927_/X _09928_/X _09930_/X vssd1 vssd1 vccd1 vccd1 _09932_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_217_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09862_ _09862_/A _09862_/B vssd1 vssd1 vccd1 vccd1 _09939_/A sky130_fd_sc_hd__nor2_8
XTAP_641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09793_ _09805_/A _09793_/B vssd1 vssd1 vccd1 vccd1 _09793_/X sky130_fd_sc_hd__or2_1
XTAP_696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_1295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_226_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_146_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09227_ _09227_/A _09227_/B _09227_/C _09227_/D vssd1 vssd1 vccd1 vccd1 _09238_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_10_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09158_ _18632_/Q _18631_/Q _18630_/Q vssd1 vssd1 vccd1 vccd1 _09160_/C sky130_fd_sc_hd__or3_4
XFILLER_177_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_182_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09089_ _18797_/Q _18796_/Q _18795_/Q vssd1 vssd1 vccd1 vccd1 _09093_/A sky130_fd_sc_hd__or3_4
XFILLER_163_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_1299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_218_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11120_ _11748_/B vssd1 vssd1 vccd1 vccd1 _13452_/A sky130_fd_sc_hd__buf_2
XFILLER_123_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11051_ _17815_/Q vssd1 vssd1 vccd1 vccd1 _11215_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_107_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_231_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10002_ _09119_/A _09114_/C _09109_/D _10350_/A _10017_/S _09709_/A vssd1 vssd1 vccd1
+ vccd1 _10002_/X sky130_fd_sc_hd__mux4_1
XFILLER_118_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14810_ _14810_/A _14814_/B vssd1 vssd1 vccd1 vccd1 _14810_/Y sky130_fd_sc_hd__nand2_1
XFILLER_76_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_218_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15790_ _18562_/Q _18526_/Q _15790_/S vssd1 vssd1 vccd1 vccd1 _15790_/X sky130_fd_sc_hd__mux2_1
XTAP_4455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14741_ _18311_/Q _18275_/Q _14756_/S vssd1 vssd1 vccd1 vccd1 _14741_/X sky130_fd_sc_hd__mux2_1
XTAP_4499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11953_ _11932_/A _11976_/A _12021_/A vssd1 vssd1 vccd1 vccd1 _11961_/B sky130_fd_sc_hd__a21oi_1
XFILLER_91_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_218_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17460_ _17493_/A _17460_/B _17460_/C vssd1 vssd1 vccd1 vccd1 _17460_/X sky130_fd_sc_hd__or3_1
X_10904_ _09376_/C _09381_/B _09386_/D _09381_/D _12089_/A _12092_/A vssd1 vssd1 vccd1
+ vccd1 _10904_/X sky130_fd_sc_hd__mux4_1
XTAP_3798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14672_ _14672_/A _14685_/B vssd1 vssd1 vccd1 vccd1 _16945_/A sky130_fd_sc_hd__or2_4
XFILLER_32_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11884_ _18159_/Q _11852_/X _11870_/Y vssd1 vssd1 vccd1 vccd1 _11885_/B sky130_fd_sc_hd__a21oi_1
XFILLER_205_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16411_ _16434_/A _16703_/B _16422_/C vssd1 vssd1 vccd1 vccd1 _16411_/X sky130_fd_sc_hd__or3_1
XFILLER_189_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13623_ _13623_/A vssd1 vssd1 vccd1 vccd1 _13624_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_73_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17391_ _18946_/Q _18910_/Q _17406_/S vssd1 vssd1 vccd1 vccd1 _17391_/X sky130_fd_sc_hd__mux2_1
X_10835_ _09253_/A _09248_/C _09243_/D _09253_/D _10702_/A _10695_/X vssd1 vssd1 vccd1
+ vccd1 _10835_/X sky130_fd_sc_hd__mux4_2
XFILLER_220_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19130_ _19130_/A _09056_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[0] sky130_fd_sc_hd__ebufn_8
XFILLER_73_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16342_ _16392_/A _16342_/B vssd1 vssd1 vccd1 vccd1 _16342_/Y sky130_fd_sc_hd__nand2_1
XFILLER_197_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13554_ _13758_/A vssd1 vssd1 vccd1 vccd1 _13573_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_125_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_164_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10766_ _10766_/A _10766_/B vssd1 vssd1 vccd1 vccd1 _10773_/A sky130_fd_sc_hd__nor2_1
XFILLER_201_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_200_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12505_ _12521_/A vssd1 vssd1 vccd1 vccd1 _17519_/A sky130_fd_sc_hd__buf_2
X_16273_ _16273_/A vssd1 vssd1 vccd1 vccd1 _16354_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_157_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_199_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10697_ _09198_/B _09193_/B _09203_/C _09193_/C _10695_/X _10852_/A vssd1 vssd1 vccd1
+ vccd1 _10697_/X sky130_fd_sc_hd__mux4_1
XFILLER_12_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13485_ _13485_/A _13526_/C _13518_/A vssd1 vssd1 vccd1 vccd1 _13563_/B sky130_fd_sc_hd__or3b_4
XFILLER_157_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18012_ _18035_/CLK _18012_/D vssd1 vssd1 vccd1 vccd1 _18012_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_201_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15224_ _15283_/A vssd1 vssd1 vccd1 vccd1 _15224_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_145_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_185_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12436_ _17901_/Q _12450_/B vssd1 vssd1 vccd1 vccd1 _12437_/B sky130_fd_sc_hd__nor2_1
XFILLER_8_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15155_ _18377_/Q _15154_/B _15154_/Y _15143_/X vssd1 vssd1 vccd1 vccd1 _18377_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_154_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12367_ _17892_/Q _17891_/Q _12444_/B _12365_/X _12366_/X vssd1 vssd1 vccd1 vccd1
+ _12369_/B sky130_fd_sc_hd__o311ai_4
XFILLER_181_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14106_ _18776_/Q _14019_/A _13625_/X _18782_/Q vssd1 vssd1 vccd1 vccd1 _14106_/X
+ sky130_fd_sc_hd__a22o_1
X_11318_ _11318_/A vssd1 vssd1 vccd1 vccd1 _11622_/A sky130_fd_sc_hd__buf_2
XFILLER_10_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15086_ _15105_/A vssd1 vssd1 vccd1 vccd1 _15100_/S sky130_fd_sc_hd__clkbuf_2
X_12298_ _11323_/A _11323_/B _11346_/A vssd1 vssd1 vccd1 vccd1 _12299_/C sky130_fd_sc_hd__o21a_1
XFILLER_141_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14037_ _18314_/Q _13625_/X _13592_/X _18332_/Q _14036_/X vssd1 vssd1 vccd1 vccd1
+ _14037_/X sky130_fd_sc_hd__a221o_1
X_11249_ _17795_/Q _17796_/Q vssd1 vssd1 vccd1 vccd1 _11404_/B sky130_fd_sc_hd__or2_2
X_18914_ _18914_/CLK _18914_/D vssd1 vssd1 vccd1 vccd1 _18914_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_95_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_228_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18845_ _18845_/CLK _18845_/D vssd1 vssd1 vccd1 vccd1 _18845_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_41_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_227_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18776_ _18778_/CLK _18776_/D vssd1 vssd1 vccd1 vccd1 _18776_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_227_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15988_ _16028_/A vssd1 vssd1 vccd1 vccd1 _15988_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_94_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17727_ _17727_/A vssd1 vssd1 vccd1 vccd1 _19007_/D sky130_fd_sc_hd__clkbuf_1
X_14939_ _18360_/Q _18324_/Q _14955_/S vssd1 vssd1 vccd1 vccd1 _14939_/X sky130_fd_sc_hd__mux2_1
XFILLER_209_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_224_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17658_ _17645_/X _17649_/Y _17654_/X _17650_/Y _18977_/Q vssd1 vssd1 vccd1 vccd1
+ _17659_/B sky130_fd_sc_hd__a32o_1
XFILLER_36_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16609_ _16611_/B _16607_/X _16608_/Y _16600_/X vssd1 vssd1 vccd1 vccd1 _18721_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_211_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17589_ _17640_/A vssd1 vssd1 vccd1 vccd1 _17610_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_91_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_204_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09012_ _09016_/A vssd1 vssd1 vccd1 vccd1 _09012_/Y sky130_fd_sc_hd__inv_2
XFILLER_178_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_219_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_208_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09914_ _09376_/C _09381_/B _09386_/D _09381_/D _09909_/X _12121_/A vssd1 vssd1 vccd1
+ vccd1 _09914_/X sky130_fd_sc_hd__mux4_1
XFILLER_217_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_219_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_217_1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09845_ _18113_/Q _17782_/Q vssd1 vssd1 vccd1 vccd1 _09846_/B sky130_fd_sc_hd__or2_1
XFILLER_86_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09776_ _09774_/A _09774_/B _09919_/A vssd1 vssd1 vccd1 vccd1 _09892_/A sky130_fd_sc_hd__o21ai_4
XTAP_3006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_4_8_0_wb_clk_i clkbuf_4_9_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_4_8_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_26_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_202_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10620_ _10731_/A _10731_/B _10619_/Y vssd1 vssd1 vccd1 vccd1 _10706_/B sky130_fd_sc_hd__a21oi_4
XFILLER_169_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10551_ _09198_/B _09193_/B _10560_/S vssd1 vssd1 vccd1 vccd1 _10552_/B sky130_fd_sc_hd__mux2_1
XFILLER_122_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13270_ _18088_/Q _12718_/X _13269_/X _13074_/X vssd1 vssd1 vccd1 vccd1 _18088_/D
+ sky130_fd_sc_hd__o211a_1
X_10482_ _10468_/X _10472_/X _10481_/X _10271_/B vssd1 vssd1 vccd1 vccd1 _10482_/X
+ sky130_fd_sc_hd__o31a_1
XFILLER_211_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12221_ _12221_/A vssd1 vssd1 vccd1 vccd1 _12221_/Y sky130_fd_sc_hd__inv_2
XFILLER_191_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12152_ _12183_/B _12154_/B _12171_/C vssd1 vssd1 vccd1 vccd1 _12152_/X sky130_fd_sc_hd__or3b_1
XFILLER_162_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19104__75 vssd1 vssd1 vccd1 vccd1 _19104__75/HI _19212_/A sky130_fd_sc_hd__conb_1
XFILLER_150_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_169_wb_clk_i clkbuf_5_10_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18094_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_11103_ _17796_/Q vssd1 vssd1 vccd1 vccd1 _11466_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_81_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16960_ _17536_/A _16960_/B vssd1 vssd1 vccd1 vccd1 _16972_/B sky130_fd_sc_hd__nor2_1
X_12083_ _12083_/A _12083_/B vssd1 vssd1 vccd1 vccd1 _12084_/B sky130_fd_sc_hd__xnor2_2
XFILLER_151_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15911_ _15938_/A _15913_/B vssd1 vssd1 vccd1 vccd1 _15911_/Y sky130_fd_sc_hd__nand2_1
X_11034_ _17972_/Q _17971_/Q vssd1 vssd1 vccd1 vccd1 _11035_/B sky130_fd_sc_hd__or2_2
XFILLER_89_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16891_ _16891_/A vssd1 vssd1 vccd1 vccd1 _17323_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_209_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18630_ _18633_/CLK _18630_/D vssd1 vssd1 vccd1 vccd1 _18630_/Q sky130_fd_sc_hd__dfxtp_2
X_15842_ _15925_/A vssd1 vssd1 vccd1 vccd1 _15842_/X sky130_fd_sc_hd__clkbuf_2
XTAP_4230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18561_ _18572_/CLK _18561_/D vssd1 vssd1 vccd1 vccd1 _18561_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_4274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15773_ _15883_/A vssd1 vssd1 vccd1 vccd1 _15863_/A sky130_fd_sc_hd__clkbuf_2
XTAP_4285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12985_ _12982_/A _12952_/X _12984_/X _12964_/X vssd1 vssd1 vccd1 vccd1 _17977_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_4296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17512_ _17512_/A _17512_/B vssd1 vssd1 vccd1 vccd1 _17512_/Y sky130_fd_sc_hd__nand2_1
XFILLER_206_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14724_ _14729_/B _14722_/X _14723_/X _14716_/X vssd1 vssd1 vccd1 vccd1 _18270_/D
+ sky130_fd_sc_hd__o211a_1
X_18492_ _18497_/CLK _18492_/D vssd1 vssd1 vccd1 vccd1 _18492_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_217_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11936_ _11975_/A _11942_/A vssd1 vssd1 vccd1 vccd1 _11984_/B sky130_fd_sc_hd__xor2_2
XFILLER_220_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17443_ _18959_/Q _18923_/Q _17447_/S vssd1 vssd1 vccd1 vccd1 _17443_/X sky130_fd_sc_hd__mux2_1
XTAP_2872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14655_ _18255_/Q _14658_/B _14654_/X _14647_/X vssd1 vssd1 vccd1 vccd1 _18255_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_127_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11867_ _11867_/A vssd1 vssd1 vccd1 vccd1 _11867_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_221_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13606_ _18837_/Q _13837_/A _13531_/A _18831_/Q vssd1 vssd1 vccd1 vccd1 _13606_/X
+ sky130_fd_sc_hd__a22o_1
X_17374_ _17514_/A _17397_/B vssd1 vssd1 vccd1 vccd1 _17383_/B sky130_fd_sc_hd__nor2_2
X_10818_ _10818_/A _10818_/B _10818_/C vssd1 vssd1 vccd1 vccd1 _10819_/D sky130_fd_sc_hd__or3_1
XFILLER_159_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14586_ _14604_/A _14589_/B vssd1 vssd1 vccd1 vccd1 _14586_/Y sky130_fd_sc_hd__nand2_1
XFILLER_20_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11798_ _11794_/X _11796_/X _11784_/X _11763_/X _11797_/Y vssd1 vssd1 vccd1 vccd1
+ _11798_/X sky130_fd_sc_hd__o221a_1
XFILLER_201_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16325_ _16325_/A _16329_/B vssd1 vssd1 vccd1 vccd1 _16325_/Y sky130_fd_sc_hd__nand2_1
XFILLER_186_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_229_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13537_ _13537_/A vssd1 vssd1 vccd1 vccd1 _13538_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_13_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_186_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10749_ _10616_/Y _10740_/X _10744_/X _10748_/X vssd1 vssd1 vccd1 vccd1 _10749_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_199_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16256_ _16268_/A _16256_/B vssd1 vssd1 vccd1 vccd1 _16256_/Y sky130_fd_sc_hd__nand2_1
XFILLER_173_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13468_ _17842_/Q _13459_/X _12184_/X vssd1 vssd1 vccd1 vccd1 _18157_/D sky130_fd_sc_hd__o21a_1
XFILLER_51_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15207_ _15207_/A vssd1 vssd1 vccd1 vccd1 _15283_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_127_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12419_ _12419_/A vssd1 vssd1 vccd1 vccd1 _12439_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_16187_ _18656_/Q _18620_/Q _16192_/S vssd1 vssd1 vccd1 vccd1 _16187_/X sky130_fd_sc_hd__mux2_1
XFILLER_57_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13399_ _18125_/Q _13398_/Y _13405_/B _11026_/X _11045_/X vssd1 vssd1 vccd1 vccd1
+ _18125_/D sky130_fd_sc_hd__o2111a_1
XFILLER_138_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15138_ _18409_/Q _18373_/Q _15141_/S vssd1 vssd1 vccd1 vccd1 _15138_/X sky130_fd_sc_hd__mux2_1
XFILLER_126_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15069_ _15115_/A _15072_/B vssd1 vssd1 vccd1 vccd1 _15069_/Y sky130_fd_sc_hd__nand2_1
XFILLER_141_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09630_ _09684_/A _09630_/B vssd1 vssd1 vccd1 vccd1 _09669_/B sky130_fd_sc_hd__xor2_4
X_18828_ _18849_/CLK _18828_/D vssd1 vssd1 vccd1 vccd1 _18828_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_28_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09561_ _18103_/Q vssd1 vssd1 vccd1 vccd1 _09580_/A sky130_fd_sc_hd__buf_2
X_18759_ _18759_/CLK _18759_/D vssd1 vssd1 vccd1 vccd1 _18759_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_55_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_224_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09492_ _18131_/Q _13357_/B vssd1 vssd1 vccd1 vccd1 _14383_/A sky130_fd_sc_hd__and2_1
XFILLER_224_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_224_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_176_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_178_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_219_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_219_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_219_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_215_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_219_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_219_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09828_ _10623_/A _09828_/B vssd1 vssd1 vccd1 vccd1 _09828_/X sky130_fd_sc_hd__and2_1
XFILLER_98_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_228_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_228_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09759_ _09760_/A _09760_/B vssd1 vssd1 vccd1 vccd1 _09784_/B sky130_fd_sc_hd__xnor2_1
XFILLER_185_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12770_ _18993_/Q vssd1 vssd1 vccd1 vccd1 _12770_/Y sky130_fd_sc_hd__inv_2
XTAP_1401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_230_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11721_ _17914_/Q vssd1 vssd1 vccd1 vccd1 _11727_/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14440_ _17564_/A _14440_/B vssd1 vssd1 vccd1 vccd1 _14441_/A sky130_fd_sc_hd__and2_1
X_11652_ _11652_/A _11652_/B vssd1 vssd1 vccd1 vccd1 _11653_/B sky130_fd_sc_hd__nor2_2
XTAP_1489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10603_ _09712_/X _09713_/X _09714_/X _09715_/X _09959_/A _10274_/S vssd1 vssd1 vccd1
+ vccd1 _10603_/X sky130_fd_sc_hd__mux4_2
XFILLER_211_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14371_ _18185_/Q _14381_/A _18186_/Q vssd1 vssd1 vccd1 vccd1 _14371_/X sky130_fd_sc_hd__o21a_1
XFILLER_183_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11583_ _11653_/A _11795_/B vssd1 vssd1 vccd1 vccd1 _11784_/B sky130_fd_sc_hd__nand2_1
XFILLER_156_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16110_ _16109_/B _16108_/X _16109_/Y _16097_/X vssd1 vssd1 vccd1 vccd1 _18602_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_11_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13322_ _18092_/Q _13322_/B vssd1 vssd1 vccd1 vccd1 _13322_/Y sky130_fd_sc_hd__nand2_1
XFILLER_11_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17090_ _18872_/Q _18836_/Q _17094_/S vssd1 vssd1 vccd1 vccd1 _17090_/X sky130_fd_sc_hd__mux2_1
X_10534_ _10547_/A _10271_/B _10526_/X _10532_/X _10533_/Y vssd1 vssd1 vccd1 vccd1
+ _10534_/X sky130_fd_sc_hd__a32o_1
XFILLER_156_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16041_ _16041_/A _16041_/B vssd1 vssd1 vccd1 vccd1 _16051_/B sky130_fd_sc_hd__nor2_2
X_13253_ _13255_/A _18081_/Q vssd1 vssd1 vccd1 vccd1 _13254_/A sky130_fd_sc_hd__and2_1
XFILLER_108_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10465_ _09287_/B _09282_/C _09282_/A _09287_/C _10464_/X _10411_/A vssd1 vssd1 vccd1
+ vccd1 _10465_/X sky130_fd_sc_hd__mux4_1
XFILLER_182_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12204_ _17853_/Q _17850_/Q _12201_/X vssd1 vssd1 vccd1 vccd1 _12210_/B sky130_fd_sc_hd__a21oi_1
XFILLER_135_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13184_ _13186_/A _18050_/Q vssd1 vssd1 vccd1 vccd1 _13185_/A sky130_fd_sc_hd__and2_1
X_10396_ _09270_/A _10813_/A _09265_/C _09265_/A _10349_/S _09969_/A vssd1 vssd1 vccd1
+ vccd1 _10396_/X sky130_fd_sc_hd__mux4_1
XFILLER_151_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12135_ _11920_/Y _12040_/X _12054_/X _12105_/X _12134_/X vssd1 vssd1 vccd1 vccd1
+ _12144_/S sky130_fd_sc_hd__o311a_4
X_17992_ _18151_/CLK _17992_/D vssd1 vssd1 vccd1 vccd1 _17992_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_96_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16943_ _16957_/A _16943_/B vssd1 vssd1 vccd1 vccd1 _16943_/Y sky130_fd_sc_hd__nand2_1
XFILLER_150_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12066_ _12066_/A _13420_/A vssd1 vssd1 vccd1 vccd1 _12066_/Y sky130_fd_sc_hd__nand2_1
XFILLER_133_1243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11017_ _11017_/A vssd1 vssd1 vccd1 vccd1 _18114_/D sky130_fd_sc_hd__clkbuf_1
X_16874_ _16884_/A _16874_/B vssd1 vssd1 vccd1 vccd1 _16874_/Y sky130_fd_sc_hd__nand2_1
XFILLER_133_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15825_ _15885_/A vssd1 vssd1 vccd1 vccd1 _15873_/A sky130_fd_sc_hd__buf_2
X_18613_ _18614_/CLK _18613_/D vssd1 vssd1 vccd1 vccd1 _18613_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_93_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_225_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_206_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18544_ _18582_/CLK _18544_/D vssd1 vssd1 vccd1 vccd1 _18544_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_3370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15756_ _18176_/Q _18175_/Q _15607_/C vssd1 vssd1 vccd1 vccd1 _17549_/A sky130_fd_sc_hd__or3b_4
XFILLER_18_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12968_ _12969_/A _12969_/B _12969_/C vssd1 vssd1 vccd1 vccd1 _12970_/A sky130_fd_sc_hd__o21a_1
Xclkbuf_leaf_66_wb_clk_i clkbuf_5_21_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18686_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_3381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14707_ _14772_/A vssd1 vssd1 vccd1 vccd1 _14843_/C sky130_fd_sc_hd__buf_2
X_18475_ _18506_/CLK _18475_/D vssd1 vssd1 vccd1 vccd1 _18475_/Q sky130_fd_sc_hd__dfxtp_2
X_11919_ _11919_/A _11919_/B vssd1 vssd1 vccd1 vccd1 _11920_/B sky130_fd_sc_hd__xnor2_4
XFILLER_221_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_206_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15687_ _15869_/A vssd1 vssd1 vccd1 vccd1 _15734_/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12899_ _17963_/Q _12899_/B vssd1 vssd1 vccd1 vccd1 _12904_/C sky130_fd_sc_hd__and2_1
XFILLER_209_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17426_ _17432_/B _17424_/X _17425_/X _17421_/X vssd1 vssd1 vccd1 vccd1 _18918_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_178_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14638_ _16905_/A vssd1 vssd1 vccd1 vccd1 _15229_/A sky130_fd_sc_hd__buf_8
XFILLER_220_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_220_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17357_ _17392_/A _17360_/B vssd1 vssd1 vccd1 vccd1 _17357_/Y sky130_fd_sc_hd__nand2_1
X_14569_ _16839_/A vssd1 vssd1 vccd1 vccd1 _15175_/B sky130_fd_sc_hd__buf_8
XFILLER_20_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_119_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16308_ _16327_/A vssd1 vssd1 vccd1 vccd1 _16324_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_9_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_201_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17288_ _17291_/B _17285_/X _17287_/Y _17283_/X vssd1 vssd1 vccd1 vccd1 _18883_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_88_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19027_ _19027_/CLK _19027_/D vssd1 vssd1 vccd1 vccd1 _19027_/Q sky130_fd_sc_hd__dfxtp_2
X_16239_ _18667_/Q _18631_/Q _16250_/S vssd1 vssd1 vccd1 vccd1 _16239_/X sky130_fd_sc_hd__mux2_1
XFILLER_47_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_216_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08992_ _08998_/A vssd1 vssd1 vccd1 vccd1 _08997_/A sky130_fd_sc_hd__buf_12
XFILLER_134_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_1351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19095__66 vssd1 vssd1 vccd1 vccd1 _19095__66/HI _19203_/A sky130_fd_sc_hd__conb_1
XFILLER_151_1310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_1354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_228_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09613_ _18126_/Q vssd1 vssd1 vccd1 vccd1 _09822_/A sky130_fd_sc_hd__buf_2
XFILLER_228_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09544_ _18103_/Q vssd1 vssd1 vccd1 vccd1 _09544_/Y sky130_fd_sc_hd__inv_2
XFILLER_3_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_225_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_212_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_224_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09475_ _09475_/A _09475_/B vssd1 vssd1 vccd1 vccd1 _09482_/B sky130_fd_sc_hd__or2_2
XFILLER_52_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_212_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_196_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_221_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_192_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_106_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10250_ _10253_/A _13348_/A _10829_/A vssd1 vssd1 vccd1 vccd1 _10250_/X sky130_fd_sc_hd__or3_1
XFILLER_117_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10181_ _10181_/A _10440_/B vssd1 vssd1 vccd1 vccd1 _10438_/A sky130_fd_sc_hd__xnor2_2
XFILLER_191_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13940_ _13940_/A vssd1 vssd1 vccd1 vccd1 _13940_/X sky130_fd_sc_hd__buf_6
XFILLER_8_1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13871_ _18451_/Q _14019_/A _13625_/X _18457_/Q _13870_/X vssd1 vssd1 vccd1 vccd1
+ _13871_/X sky130_fd_sc_hd__a221o_1
XFILLER_19_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15610_ _16055_/A _15748_/C vssd1 vssd1 vccd1 vccd1 _15618_/B sky130_fd_sc_hd__nor2_2
XFILLER_189_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12822_ _12570_/B _12816_/X _12818_/X _12821_/Y vssd1 vssd1 vccd1 vccd1 _12822_/X
+ sky130_fd_sc_hd__a211o_1
X_16590_ _18716_/Q _16589_/B _16589_/Y _16581_/X vssd1 vssd1 vccd1 vccd1 _18716_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_90_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_215_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15541_ _15546_/B _15539_/X _15540_/X _15536_/X vssd1 vssd1 vccd1 vccd1 _18465_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_188_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_231_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_203_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12753_ _18013_/Q _18012_/Q _18015_/Q _18014_/Q vssd1 vssd1 vccd1 vccd1 _12754_/D
+ sky130_fd_sc_hd__and4_1
XFILLER_43_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_5_17_0_wb_clk_i clkbuf_4_8_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18759_/CLK
+ sky130_fd_sc_hd__clkbuf_2
XTAP_1242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18260_ _18266_/CLK _18260_/D vssd1 vssd1 vccd1 vccd1 _18260_/Q sky130_fd_sc_hd__dfxtp_1
X_11704_ _11704_/A _11704_/B _11704_/C _11619_/X vssd1 vssd1 vccd1 vccd1 _11705_/C
+ sky130_fd_sc_hd__or4b_1
XFILLER_15_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_231_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_187_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15472_ _18448_/Q _15473_/B _15471_/Y _15452_/X vssd1 vssd1 vccd1 vccd1 _18448_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_1275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12684_ _17936_/Q vssd1 vssd1 vccd1 vccd1 _12697_/B sky130_fd_sc_hd__clkinv_2
XTAP_1286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17211_ _17213_/B _17209_/X _17210_/Y _17197_/X vssd1 vssd1 vccd1 vccd1 _18865_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_230_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14423_ _14423_/A vssd1 vssd1 vccd1 vccd1 _14423_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_202_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11635_ _11635_/A _11757_/A _11635_/C vssd1 vssd1 vccd1 vccd1 _11635_/X sky130_fd_sc_hd__or3_2
X_18191_ _18191_/CLK _18191_/D vssd1 vssd1 vccd1 vccd1 _18191_/Q sky130_fd_sc_hd__dfxtp_1
X_17142_ _18884_/Q _18848_/Q _17151_/S vssd1 vssd1 vccd1 vccd1 _17142_/X sky130_fd_sc_hd__mux2_1
X_14354_ _14584_/A vssd1 vssd1 vccd1 vccd1 _14354_/X sky130_fd_sc_hd__buf_4
XFILLER_11_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11566_ _11549_/X _11563_/C _11565_/X vssd1 vssd1 vccd1 vccd1 _11566_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_183_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_184_wb_clk_i clkbuf_5_8_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _19019_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_13305_ _18081_/Q _18080_/Q _18083_/Q _18082_/Q vssd1 vssd1 vccd1 vccd1 _13310_/B
+ sky130_fd_sc_hd__or4_1
X_17073_ _17080_/B _17071_/X _17072_/X _17057_/X vssd1 vssd1 vccd1 vccd1 _18831_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_116_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10517_ _10439_/X _10516_/Y _10939_/A vssd1 vssd1 vccd1 vccd1 _13411_/B sky130_fd_sc_hd__a21oi_1
XFILLER_196_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14285_ _15607_/B vssd1 vssd1 vccd1 vccd1 _15145_/B sky130_fd_sc_hd__buf_4
XFILLER_157_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11497_ _11654_/C _11497_/B vssd1 vssd1 vccd1 vccd1 _11499_/B sky130_fd_sc_hd__or2_1
XFILLER_109_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_113_wb_clk_i clkbuf_5_31_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18497_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_16024_ _16062_/A _16027_/B vssd1 vssd1 vccd1 vccd1 _16024_/Y sky130_fd_sc_hd__nand2_1
XFILLER_171_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13236_ _13244_/A _18073_/Q vssd1 vssd1 vccd1 vccd1 _13237_/A sky130_fd_sc_hd__and2_1
XFILLER_100_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10448_ _10560_/S vssd1 vssd1 vccd1 vccd1 _10550_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_108_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13167_ _13175_/A _18042_/Q vssd1 vssd1 vccd1 vccd1 _13168_/A sky130_fd_sc_hd__and2_1
XFILLER_69_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10379_ _09332_/B _09327_/B _09337_/C _09327_/C _09945_/X _09905_/X vssd1 vssd1 vccd1
+ vccd1 _10379_/X sky130_fd_sc_hd__mux4_2
XFILLER_83_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12118_ _12118_/A _12118_/B vssd1 vssd1 vccd1 vccd1 _12119_/B sky130_fd_sc_hd__xnor2_2
X_13098_ _13142_/A vssd1 vssd1 vccd1 vccd1 _13107_/A sky130_fd_sc_hd__clkbuf_1
X_17975_ _18108_/CLK _17975_/D vssd1 vssd1 vccd1 vccd1 _17975_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_97_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16926_ _16954_/A _16930_/B vssd1 vssd1 vccd1 vccd1 _16926_/Y sky130_fd_sc_hd__nand2_1
X_12049_ _12049_/A _12049_/B vssd1 vssd1 vccd1 vccd1 _12055_/B sky130_fd_sc_hd__and2_4
XFILLER_111_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16857_ _16882_/A _16860_/B vssd1 vssd1 vccd1 vccd1 _16857_/Y sky130_fd_sc_hd__nand2_1
XFILLER_225_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19038__9 vssd1 vssd1 vccd1 vccd1 _19038__9/HI _19132_/A sky130_fd_sc_hd__conb_1
X_15808_ _15962_/A _15844_/B vssd1 vssd1 vccd1 vccd1 _15818_/B sky130_fd_sc_hd__nor2_1
XFILLER_168_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16788_ _18802_/Q _18766_/Q _16802_/S vssd1 vssd1 vccd1 vccd1 _16788_/X sky130_fd_sc_hd__mux2_1
XFILLER_81_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_1333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18527_ _18563_/CLK _18527_/D vssd1 vssd1 vccd1 vccd1 _18527_/Q sky130_fd_sc_hd__dfxtp_4
X_15739_ _15739_/A vssd1 vssd1 vccd1 vccd1 _15823_/A sky130_fd_sc_hd__buf_2
XFILLER_45_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_1306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09260_ _09260_/A _09260_/B _10317_/A _09260_/D vssd1 vssd1 vccd1 vccd1 _09271_/A
+ sky130_fd_sc_hd__and4_1
X_18458_ _18458_/CLK _18458_/D vssd1 vssd1 vccd1 vccd1 _18458_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_209_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_181_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_221_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09191_ _18575_/Q _18574_/Q _18573_/Q vssd1 vssd1 vccd1 vccd1 _09193_/C sky130_fd_sc_hd__or3_4
XFILLER_60_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17409_ _17408_/B _17406_/X _17408_/Y _17400_/X vssd1 vssd1 vccd1 vccd1 _18914_/D
+ sky130_fd_sc_hd__o211a_1
X_18389_ _18398_/CLK _18389_/D vssd1 vssd1 vccd1 vccd1 _18389_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_187_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_216_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08975_ _08979_/A vssd1 vssd1 vccd1 vccd1 _08975_/Y sky130_fd_sc_hd__inv_2
XFILLER_25_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_225_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09527_ _18112_/Q vssd1 vssd1 vccd1 vccd1 _10113_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_227_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09458_ _09458_/A vssd1 vssd1 vccd1 vccd1 _18131_/D sky130_fd_sc_hd__clkbuf_1
XPHY_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_223_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_212_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_212_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09389_ _18347_/Q _18346_/Q _18345_/Q vssd1 vssd1 vccd1 vccd1 _09392_/B sky130_fd_sc_hd__or3_2
XFILLER_61_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11420_ _12329_/A _12316_/B _11338_/A _11419_/X vssd1 vssd1 vccd1 vccd1 _11420_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_32_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_184_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_197_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11351_ _13447_/A _11748_/B _11495_/D vssd1 vssd1 vccd1 vccd1 _11593_/B sky130_fd_sc_hd__nand3b_4
XFILLER_192_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_165_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10302_ _09186_/A _09181_/A _09181_/D _09176_/D _09947_/A _10599_/S vssd1 vssd1 vccd1
+ vccd1 _10302_/X sky130_fd_sc_hd__mux4_2
XFILLER_158_1349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14070_ _18827_/Q _13596_/X _13630_/X _18809_/Q vssd1 vssd1 vccd1 vccd1 _14070_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_125_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11282_ _11905_/A _11282_/B _11812_/B _11281_/X vssd1 vssd1 vccd1 vccd1 _11869_/A
+ sky130_fd_sc_hd__nor4b_2
XFILLER_134_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13021_ _17984_/Q _13036_/B vssd1 vssd1 vccd1 vccd1 _13021_/X sky130_fd_sc_hd__or2_1
XFILLER_106_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10233_ _10521_/A vssd1 vssd1 vccd1 vccd1 _10542_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_10_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10164_ _17982_/Q vssd1 vssd1 vccd1 vccd1 _13009_/A sky130_fd_sc_hd__buf_4
XFILLER_120_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14972_ _14971_/B _14970_/X _14971_/Y _14961_/X vssd1 vssd1 vccd1 vccd1 _18332_/D
+ sky130_fd_sc_hd__o211a_1
X_17760_ _17764_/A _19024_/Q vssd1 vssd1 vccd1 vccd1 _17761_/A sky130_fd_sc_hd__and2_1
X_10095_ _09253_/A _09248_/C _09243_/D _09253_/D _09995_/A _09708_/A vssd1 vssd1 vccd1
+ vccd1 _10095_/X sky130_fd_sc_hd__mux4_1
XFILLER_59_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13923_ _13916_/X _13922_/X _13710_/Y vssd1 vssd1 vccd1 vccd1 _13923_/X sky130_fd_sc_hd__o21a_2
X_16711_ _16832_/A vssd1 vssd1 vccd1 vccd1 _16755_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_47_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17691_ _17691_/A vssd1 vssd1 vccd1 vccd1 _18984_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_19_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16642_ _18766_/Q _18730_/Q _16657_/S vssd1 vssd1 vccd1 vccd1 _16642_/X sky130_fd_sc_hd__mux2_1
XFILLER_90_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13854_ _18706_/Q _13577_/X _13850_/X _13853_/X vssd1 vssd1 vccd1 vccd1 _13854_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_207_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_223_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12805_ _12609_/B _12871_/A _12802_/Y _12627_/B _12804_/X vssd1 vssd1 vccd1 vccd1
+ _12813_/B sky130_fd_sc_hd__o221ai_1
XFILLER_76_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_204_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16573_ _16575_/B _16571_/X _16572_/Y _16559_/X vssd1 vssd1 vccd1 vccd1 _18712_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_16_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13785_ _13785_/A vssd1 vssd1 vccd1 vccd1 _13785_/X sky130_fd_sc_hd__buf_8
XFILLER_90_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10997_ _17819_/Q vssd1 vssd1 vccd1 vccd1 _11232_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_188_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15524_ _15582_/A vssd1 vssd1 vccd1 vccd1 _15570_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_203_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18312_ _18312_/CLK _18312_/D vssd1 vssd1 vccd1 vccd1 _18312_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_206_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12736_ _12736_/A _12736_/B _12736_/C vssd1 vssd1 vccd1 vccd1 _12743_/B sky130_fd_sc_hd__and3_1
XTAP_1061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18243_ _18244_/CLK _18243_/D vssd1 vssd1 vccd1 vccd1 _18243_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15455_ _15578_/A vssd1 vssd1 vccd1 vccd1 _15508_/A sky130_fd_sc_hd__buf_2
XFILLER_163_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12667_ _12708_/A vssd1 vssd1 vccd1 vccd1 _12667_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_175_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14406_ _14404_/X _09495_/B _14405_/X vssd1 vssd1 vccd1 vccd1 _14406_/X sky130_fd_sc_hd__a21o_1
XFILLER_15_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11618_ _11603_/Y _11616_/Y _11617_/X vssd1 vssd1 vccd1 vccd1 _11618_/Y sky130_fd_sc_hd__a21oi_1
X_18174_ _18182_/CLK _18174_/D vssd1 vssd1 vccd1 vccd1 _18174_/Q sky130_fd_sc_hd__dfxtp_1
X_15386_ _15442_/A _15390_/B vssd1 vssd1 vccd1 vccd1 _15386_/Y sky130_fd_sc_hd__nand2_1
XFILLER_156_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12598_ _12598_/A _12598_/B vssd1 vssd1 vccd1 vccd1 _12600_/B sky130_fd_sc_hd__nor2_1
XFILLER_50_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17125_ _17136_/A _17415_/B _17173_/C vssd1 vssd1 vccd1 vccd1 _17125_/X sky130_fd_sc_hd__or3_1
XFILLER_7_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14337_ _14349_/A _14333_/X _14334_/Y _14336_/X vssd1 vssd1 vccd1 vccd1 _14337_/X
+ sky130_fd_sc_hd__o31a_1
XFILLER_102_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11549_ _19032_/Q vssd1 vssd1 vccd1 vccd1 _11549_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_116_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_183_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17056_ _17091_/A _17056_/B vssd1 vssd1 vccd1 vccd1 _17056_/Y sky130_fd_sc_hd__nand2_1
X_14268_ _14267_/A _14266_/Y _14267_/Y _13409_/X vssd1 vssd1 vccd1 vccd1 _14268_/X
+ sky130_fd_sc_hd__o211a_1
X_16007_ _16043_/A _16007_/B _16021_/C vssd1 vssd1 vccd1 vccd1 _16007_/X sky130_fd_sc_hd__or3_1
X_13219_ _13219_/A vssd1 vssd1 vccd1 vccd1 _18064_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_143_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14199_ _14199_/A _14349_/B vssd1 vssd1 vccd1 vccd1 _14300_/A sky130_fd_sc_hd__nor2_1
XFILLER_135_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_1176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_4_10_0_wb_clk_i clkbuf_3_5_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_5_21_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_170_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19065__36 vssd1 vssd1 vccd1 vccd1 _19065__36/HI _19159_/A sky130_fd_sc_hd__conb_1
XFILLER_39_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17958_ _17959_/CLK _17958_/D vssd1 vssd1 vccd1 vccd1 _17958_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_81_wb_clk_i clkbuf_5_23_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18571_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_39_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16909_ _16909_/A vssd1 vssd1 vccd1 vccd1 _17493_/B sky130_fd_sc_hd__buf_6
X_17889_ _17890_/CLK _17889_/D vssd1 vssd1 vccd1 vccd1 _17889_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_226_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_213_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_198_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_111_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09312_ _18476_/Q _18475_/Q _18474_/Q vssd1 vssd1 vccd1 vccd1 _09314_/C sky130_fd_sc_hd__or3_4
XFILLER_0_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_221_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_222_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09243_ _09243_/A _09243_/B _09243_/C _09243_/D vssd1 vssd1 vccd1 vccd1 _09254_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_181_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09174_ _18617_/Q _18616_/Q _18615_/Q vssd1 vssd1 vccd1 vccd1 _09176_/C sky130_fd_sc_hd__or3_4
XFILLER_159_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_222_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_227_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_227_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08958_ _08960_/A vssd1 vssd1 vccd1 vccd1 _08958_/Y sky130_fd_sc_hd__inv_2
XTAP_5349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_217_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10920_ _11925_/A _10920_/B vssd1 vssd1 vccd1 vccd1 _10920_/X sky130_fd_sc_hd__and2_1
XTAP_3958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_205_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10851_ _10851_/A vssd1 vssd1 vccd1 vccd1 _14206_/A sky130_fd_sc_hd__buf_4
XFILLER_147_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_112_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_1331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_198_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13570_ _18669_/Q _13546_/X _13556_/X _13569_/X vssd1 vssd1 vccd1 vccd1 _13570_/X
+ sky130_fd_sc_hd__a211o_1
XPHY_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_227_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10782_ _10782_/A _10813_/B vssd1 vssd1 vccd1 vccd1 _10782_/X sky130_fd_sc_hd__or2_1
XFILLER_25_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12521_ _12521_/A _12528_/C vssd1 vssd1 vccd1 vccd1 _12522_/A sky130_fd_sc_hd__or2b_2
XPHY_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_227_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15240_ _15239_/B _15238_/X _15239_/Y _15224_/X vssd1 vssd1 vccd1 vccd1 _18398_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_12_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12452_ _12452_/A _12452_/B _12452_/C vssd1 vssd1 vccd1 vccd1 _12454_/B sky130_fd_sc_hd__nand3_1
XFILLER_173_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_200_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11403_ _11403_/A _11497_/B vssd1 vssd1 vccd1 vccd1 _11412_/A sky130_fd_sc_hd__nor2_1
X_15171_ _15211_/A vssd1 vssd1 vccd1 vccd1 _15229_/B sky130_fd_sc_hd__buf_2
XFILLER_153_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12383_ _12384_/B _12384_/C _17895_/Q vssd1 vssd1 vccd1 vccd1 _12397_/A sky130_fd_sc_hd__o21a_1
XFILLER_181_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14122_ _18896_/Q _13568_/X _13842_/X _18890_/Q _14121_/X vssd1 vssd1 vccd1 vccd1
+ _14122_/X sky130_fd_sc_hd__a221o_1
XFILLER_153_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11334_ _11334_/A _11334_/B _11336_/A _11336_/B vssd1 vssd1 vccd1 vccd1 _11334_/X
+ sky130_fd_sc_hd__and4_1
XFILLER_126_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_1321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14053_ _18488_/Q _13507_/A _14030_/A _18512_/Q vssd1 vssd1 vccd1 vccd1 _14053_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_84_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18930_ _18931_/CLK _18930_/D vssd1 vssd1 vccd1 vccd1 _18930_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_180_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11265_ _11748_/B _11259_/Y _11264_/Y _11780_/A vssd1 vssd1 vccd1 vccd1 _11265_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_79_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13004_ _13005_/A _13005_/B vssd1 vssd1 vccd1 vccd1 _13004_/X sky130_fd_sc_hd__or2_1
X_10216_ _10440_/A _10227_/B vssd1 vssd1 vccd1 vccd1 _10232_/A sky130_fd_sc_hd__nor2_2
X_18861_ _18862_/CLK _18861_/D vssd1 vssd1 vccd1 vccd1 _18861_/Q sky130_fd_sc_hd__dfxtp_2
X_11196_ _17811_/Q _11196_/B _17809_/Q _11196_/D vssd1 vssd1 vccd1 vccd1 _11205_/C
+ sky130_fd_sc_hd__and4_1
XFILLER_79_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17812_ _18989_/CLK _17812_/D vssd1 vssd1 vccd1 vccd1 _17812_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_67_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10147_ _10147_/A _10147_/B vssd1 vssd1 vccd1 vccd1 _10175_/B sky130_fd_sc_hd__nor2_2
XFILLER_79_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18792_ _18812_/CLK _18792_/D vssd1 vssd1 vccd1 vccd1 _18792_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_5850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14955_ _18364_/Q _18328_/Q _14955_/S vssd1 vssd1 vccd1 vccd1 _14955_/X sky130_fd_sc_hd__mux2_1
XFILLER_134_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17743_ _17745_/A _19016_/Q vssd1 vssd1 vccd1 vccd1 _17744_/A sky130_fd_sc_hd__and2_1
X_10078_ _09093_/A _09093_/B _09098_/C _09103_/B _09703_/A _09689_/X vssd1 vssd1 vccd1
+ vccd1 _10078_/X sky130_fd_sc_hd__mux4_2
XFILLER_130_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13906_ _18877_/Q _13906_/B vssd1 vssd1 vccd1 vccd1 _13906_/X sky130_fd_sc_hd__and2_1
X_14886_ _14890_/B _14883_/X _14885_/Y _14881_/X vssd1 vssd1 vccd1 vccd1 _18310_/D
+ sky130_fd_sc_hd__o211a_1
X_17674_ _17674_/A _17687_/B vssd1 vssd1 vccd1 vccd1 _17674_/Y sky130_fd_sc_hd__nor2_1
XFILLER_208_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINSDIODE2_202 _14504_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16625_ _16771_/A _16650_/B vssd1 vssd1 vccd1 vccd1 _16634_/B sky130_fd_sc_hd__nor2_1
X_13837_ _13837_/A vssd1 vssd1 vccd1 vccd1 _13838_/A sky130_fd_sc_hd__buf_4
XINSDIODE2_213 _13630_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_224 _15150_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINSDIODE2_235 _16666_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_223_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_204_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_246 _17549_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16556_ _16562_/B _16554_/X _16555_/X _16539_/X vssd1 vssd1 vccd1 vccd1 _18708_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_189_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XINSDIODE2_257 _13575_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13768_ _18513_/Q _13738_/X _13765_/X _13767_/X vssd1 vssd1 vccd1 vccd1 _13768_/X
+ sky130_fd_sc_hd__a211o_1
XINSDIODE2_268 input1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_210_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_189_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15507_ _18493_/Q _18457_/Q _15514_/S vssd1 vssd1 vccd1 vccd1 _15507_/X sky130_fd_sc_hd__mux2_1
XFILLER_176_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12719_ _17940_/Q _18000_/Q vssd1 vssd1 vccd1 vccd1 _12926_/A sky130_fd_sc_hd__and2b_1
XFILLER_91_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16487_ _16510_/A _16487_/B vssd1 vssd1 vccd1 vccd1 _16487_/Y sky130_fd_sc_hd__nand2_1
XFILLER_149_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13699_ _18768_/Q _14014_/A _14026_/A _18759_/Q vssd1 vssd1 vccd1 vccd1 _13699_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_30_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15438_ _15492_/A _16032_/B _15451_/C vssd1 vssd1 vccd1 vccd1 _15438_/X sky130_fd_sc_hd__or3_1
X_18226_ _19026_/CLK _18226_/D vssd1 vssd1 vccd1 vccd1 _18226_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_191_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_1292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15369_ _15562_/A vssd1 vssd1 vccd1 vccd1 _15423_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_18157_ _18157_/CLK _18157_/D vssd1 vssd1 vccd1 vccd1 _18157_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_129_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_2_0_1_wb_clk_i clkbuf_2_0_1_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_1_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_2
X_17108_ _18876_/Q _18840_/Q _17114_/S vssd1 vssd1 vccd1 vccd1 _17108_/X sky130_fd_sc_hd__mux2_1
X_18088_ _18088_/CLK _18088_/D vssd1 vssd1 vccd1 vccd1 _18088_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_171_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17039_ _17072_/A _17473_/B _17085_/C vssd1 vssd1 vccd1 vccd1 _17039_/X sky130_fd_sc_hd__or3_1
X_09930_ _09930_/A vssd1 vssd1 vccd1 vccd1 _09930_/X sky130_fd_sc_hd__buf_4
XFILLER_125_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09861_ _09860_/B _09860_/C _09860_/A vssd1 vssd1 vccd1 vccd1 _09862_/B sky130_fd_sc_hd__o21a_2
XFILLER_113_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_217_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_213_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09792_ _09792_/A _09792_/B vssd1 vssd1 vccd1 vccd1 _09812_/A sky130_fd_sc_hd__xnor2_2
XFILLER_218_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_148_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_93_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_214_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_216_wb_clk_i clkbuf_5_8_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17879_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_59_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_224_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_158_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09226_ _18926_/Q _18925_/Q _18924_/Q vssd1 vssd1 vccd1 vccd1 _09227_/D sky130_fd_sc_hd__or3_4
XFILLER_139_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09157_ _18647_/Q _18646_/Q _18645_/Q vssd1 vssd1 vccd1 vccd1 _09160_/B sky130_fd_sc_hd__or3_4
XFILLER_181_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_1305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09088_ _09088_/A vssd1 vssd1 vccd1 vccd1 _19182_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_108_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_122_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11050_ _17785_/Q vssd1 vssd1 vccd1 vccd1 _11333_/A sky130_fd_sc_hd__clkbuf_2
XTAP_5102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10001_ _12068_/A _09988_/X _09997_/X _10940_/A vssd1 vssd1 vccd1 vccd1 _10001_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_49_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_231_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_191_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14740_ _14812_/A vssd1 vssd1 vccd1 vccd1 _14756_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_18_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11952_ _11970_/A _11984_/B vssd1 vssd1 vccd1 vccd1 _11999_/B sky130_fd_sc_hd__nand2_1
XTAP_4489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10903_ _10899_/X _10902_/X _10903_/S vssd1 vssd1 vccd1 vccd1 _10903_/X sky130_fd_sc_hd__mux2_1
XFILLER_205_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14671_ _18260_/Q _14670_/B _14670_/Y _14668_/X vssd1 vssd1 vccd1 vccd1 _18260_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_3788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11883_ _12207_/A _11883_/B vssd1 vssd1 vccd1 vccd1 _17833_/D sky130_fd_sc_hd__nor2_1
X_16410_ _18708_/Q _18672_/Q _16421_/S vssd1 vssd1 vccd1 vccd1 _16410_/X sky130_fd_sc_hd__mux2_1
XFILLER_205_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13622_ _13667_/A vssd1 vssd1 vccd1 vccd1 _13623_/A sky130_fd_sc_hd__buf_6
XFILLER_32_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17390_ _17390_/A vssd1 vssd1 vccd1 vccd1 _17406_/S sky130_fd_sc_hd__clkbuf_2
X_10834_ _09248_/B _09243_/B _09253_/C _09243_/C _10695_/X _10648_/X vssd1 vssd1 vccd1
+ vccd1 _10834_/X sky130_fd_sc_hd__mux4_2
XFILLER_60_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_201_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_186_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16341_ _16524_/A vssd1 vssd1 vccd1 vccd1 _16392_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_164_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_186_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13553_ _13906_/B vssd1 vssd1 vccd1 vccd1 _13758_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_160_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10765_ _10824_/A _10762_/X _10764_/X _10753_/A vssd1 vssd1 vccd1 vccd1 _10766_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_160_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12504_ _18132_/Q _13357_/B vssd1 vssd1 vccd1 vccd1 _12521_/A sky130_fd_sc_hd__nand2_1
X_16272_ _16310_/A _16716_/B _16272_/C vssd1 vssd1 vccd1 vccd1 _16272_/X sky130_fd_sc_hd__or3_1
XFILLER_185_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13484_ _17849_/Q _13459_/X _12184_/X vssd1 vssd1 vccd1 vccd1 _18165_/D sky130_fd_sc_hd__o21a_1
X_10696_ _10811_/A vssd1 vssd1 vccd1 vccd1 _10852_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_199_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15223_ _15236_/A _15227_/B vssd1 vssd1 vccd1 vccd1 _15223_/Y sky130_fd_sc_hd__nand2_1
XFILLER_139_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18011_ _19004_/CLK _18011_/D vssd1 vssd1 vccd1 vccd1 _18011_/Q sky130_fd_sc_hd__dfxtp_1
X_12435_ _17901_/Q _12450_/B vssd1 vssd1 vccd1 vccd1 _12437_/A sky130_fd_sc_hd__and2_1
XFILLER_12_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_218_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15154_ _15182_/A _15154_/B vssd1 vssd1 vccd1 vccd1 _15154_/Y sky130_fd_sc_hd__nand2_1
X_12366_ _17893_/Q _12373_/A vssd1 vssd1 vccd1 vccd1 _12366_/X sky130_fd_sc_hd__or2b_1
XFILLER_153_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14105_ _18785_/Q _13858_/X _13500_/X _18800_/Q _14104_/X vssd1 vssd1 vccd1 vccd1
+ _14105_/X sky130_fd_sc_hd__a221o_1
X_11317_ _11375_/A _11340_/B vssd1 vssd1 vccd1 vccd1 _11318_/A sky130_fd_sc_hd__nand2_2
X_15085_ _15229_/A _15085_/B vssd1 vssd1 vccd1 vccd1 _15094_/B sky130_fd_sc_hd__nor2_1
XFILLER_181_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12297_ _12297_/A vssd1 vssd1 vccd1 vccd1 _17874_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_10_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14036_ _18320_/Q _13877_/A _13642_/X _18308_/Q vssd1 vssd1 vccd1 vccd1 _14036_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_141_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18913_ _18914_/CLK _18913_/D vssd1 vssd1 vccd1 vccd1 _18913_/Q sky130_fd_sc_hd__dfxtp_1
X_11248_ _13501_/A vssd1 vssd1 vccd1 vccd1 _11653_/A sky130_fd_sc_hd__buf_2
XFILLER_106_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18844_ _18845_/CLK _18844_/D vssd1 vssd1 vccd1 vccd1 _18844_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_136_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11179_ _11179_/A vssd1 vssd1 vccd1 vccd1 _17806_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_228_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_171_1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18775_ _18778_/CLK _18775_/D vssd1 vssd1 vccd1 vccd1 _18775_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_5680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15987_ _16000_/A _15991_/B vssd1 vssd1 vccd1 vccd1 _15987_/Y sky130_fd_sc_hd__nand2_1
XTAP_5691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_212_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17726_ _17734_/A _19008_/Q vssd1 vssd1 vccd1 vccd1 _17727_/A sky130_fd_sc_hd__and2_1
X_14938_ _14958_/A vssd1 vssd1 vccd1 vccd1 _14955_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_224_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_224_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17657_ _17657_/A vssd1 vssd1 vccd1 vccd1 _18976_/D sky130_fd_sc_hd__clkbuf_1
X_14869_ _14919_/A _15162_/B _14906_/C vssd1 vssd1 vccd1 vccd1 _14869_/X sky130_fd_sc_hd__or3_1
XFILLER_35_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16608_ _16631_/A _16611_/B vssd1 vssd1 vccd1 vccd1 _16608_/Y sky130_fd_sc_hd__nand2_1
XFILLER_91_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_189_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17588_ _17588_/A vssd1 vssd1 vccd1 vccd1 _18959_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_143_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16539_ _16559_/A vssd1 vssd1 vccd1 vccd1 _16539_/X sky130_fd_sc_hd__dlymetal6s2s_1
Xclkbuf_1_1_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_1_1_1_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_52_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_176_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_149_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09011_ _09029_/A vssd1 vssd1 vccd1 vccd1 _09016_/A sky130_fd_sc_hd__buf_12
X_18209_ _18209_/CLK _18209_/D vssd1 vssd1 vccd1 vccd1 _18209_/Q sky130_fd_sc_hd__dfxtp_1
X_19189_ _19189_/A _08989_/Y vssd1 vssd1 vccd1 vccd1 io_out[27] sky130_fd_sc_hd__ebufn_8
XFILLER_128_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_171_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09913_ _09959_/A vssd1 vssd1 vccd1 vccd1 _12121_/A sky130_fd_sc_hd__buf_6
XFILLER_160_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_217_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09844_ _09844_/A _17782_/Q vssd1 vssd1 vccd1 vccd1 _09846_/A sky130_fd_sc_hd__nand2_1
XFILLER_113_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09775_ _09918_/A _09918_/B vssd1 vssd1 vccd1 vccd1 _09919_/A sky130_fd_sc_hd__or2_2
XFILLER_218_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_227_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_226_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_183_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_230_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_1178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_214_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_169_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10550_ _09203_/C _09193_/C _10550_/S vssd1 vssd1 vccd1 vccd1 _10550_/X sky130_fd_sc_hd__mux2_1
XFILLER_10_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09209_ _09209_/A _09209_/B _09209_/C _10795_/A vssd1 vssd1 vccd1 vccd1 _09220_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_6_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_202_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10481_ _10474_/X _10443_/X _10477_/X _10480_/X _10547_/B vssd1 vssd1 vccd1 vccd1
+ _10481_/X sky130_fd_sc_hd__a32o_1
XFILLER_108_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12220_ _12493_/B _12358_/B _17854_/Q _12219_/X vssd1 vssd1 vccd1 vccd1 _17854_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_108_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12151_ _12151_/A _12169_/A _12169_/B vssd1 vssd1 vccd1 vccd1 _12171_/C sky130_fd_sc_hd__or3_1
XFILLER_2_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11102_ _11102_/A vssd1 vssd1 vccd1 vccd1 _17795_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_150_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12082_ _12082_/A _12082_/B vssd1 vssd1 vccd1 vccd1 _12083_/B sky130_fd_sc_hd__xnor2_1
XFILLER_89_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15910_ _18555_/Q _15913_/B _15909_/X _15901_/X vssd1 vssd1 vccd1 vccd1 _18555_/D
+ sky130_fd_sc_hd__o211a_1
X_11033_ _17970_/Q vssd1 vssd1 vccd1 vccd1 _13368_/B sky130_fd_sc_hd__buf_2
XFILLER_81_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16890_ _16936_/A _17483_/B _16936_/C vssd1 vssd1 vccd1 vccd1 _16890_/X sky130_fd_sc_hd__or3_1
XFILLER_89_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_231_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15841_ _16273_/A vssd1 vssd1 vccd1 vccd1 _15925_/A sky130_fd_sc_hd__clkbuf_2
XTAP_4220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_218_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_138_wb_clk_i clkbuf_5_27_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18356_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_4253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18560_ _18572_/CLK _18560_/D vssd1 vssd1 vccd1 vccd1 _18560_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_4264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_224_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15772_ _18143_/Q _15772_/B vssd1 vssd1 vccd1 vccd1 _15883_/A sky130_fd_sc_hd__nand2_2
XTAP_4275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12984_ _17987_/Q _12955_/X _12983_/Y _12721_/X _12949_/Y vssd1 vssd1 vccd1 vccd1
+ _12984_/X sky130_fd_sc_hd__a221o_1
XFILLER_91_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17511_ _18977_/Q _18941_/Q _17515_/S vssd1 vssd1 vccd1 vccd1 _17511_/X sky130_fd_sc_hd__mux2_1
X_14723_ _14734_/A _15162_/B _14757_/C vssd1 vssd1 vccd1 vccd1 _14723_/X sky130_fd_sc_hd__or3_1
XFILLER_45_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11935_ _11970_/A _11951_/A vssd1 vssd1 vccd1 vccd1 _11944_/A sky130_fd_sc_hd__or2_1
X_18491_ _18496_/CLK _18491_/D vssd1 vssd1 vccd1 vccd1 _18491_/Q sky130_fd_sc_hd__dfxtp_4
XTAP_3574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14654_ _14665_/A _14665_/B _15243_/B vssd1 vssd1 vccd1 vccd1 _14654_/X sky130_fd_sc_hd__or3_1
XFILLER_45_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17442_ _17444_/B _17439_/X _17440_/Y _17441_/X vssd1 vssd1 vccd1 vccd1 _18922_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_2873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11866_ _14421_/A vssd1 vssd1 vccd1 vccd1 _11879_/A sky130_fd_sc_hd__clkbuf_2
XTAP_2884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_177_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13605_ _18810_/Q _13591_/X _13592_/X _18834_/Q _13604_/X vssd1 vssd1 vccd1 vccd1
+ _13605_/X sky130_fd_sc_hd__a221o_1
XFILLER_214_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10817_ _09270_/B _09260_/B _09260_/D _10317_/A _10668_/A _10883_/B vssd1 vssd1 vccd1
+ vccd1 _10818_/C sky130_fd_sc_hd__mux4_1
X_14585_ _18240_/Q _14589_/B _14584_/X _14561_/X vssd1 vssd1 vccd1 vccd1 _18240_/D
+ sky130_fd_sc_hd__o211a_1
X_17373_ _17372_/B _17371_/X _17372_/Y _17361_/X vssd1 vssd1 vccd1 vccd1 _18905_/D
+ sky130_fd_sc_hd__o211a_1
X_11797_ _11797_/A _11797_/B vssd1 vssd1 vccd1 vccd1 _11797_/Y sky130_fd_sc_hd__nand2_1
XFILLER_60_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16324_ _18688_/Q _18652_/Q _16324_/S vssd1 vssd1 vccd1 vccd1 _16324_/X sky130_fd_sc_hd__mux2_1
X_13536_ _13706_/A vssd1 vssd1 vccd1 vccd1 _13537_/A sky130_fd_sc_hd__clkbuf_8
X_10748_ _10738_/A _10745_/X _10747_/X _10733_/A vssd1 vssd1 vccd1 vccd1 _10748_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_201_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_229_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_186_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16255_ _18671_/Q _18635_/Q _16271_/S vssd1 vssd1 vccd1 vccd1 _16255_/X sky130_fd_sc_hd__mux2_1
XFILLER_145_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13467_ _13467_/A _13467_/B vssd1 vssd1 vccd1 vccd1 _18156_/D sky130_fd_sc_hd__nor2_1
XFILLER_51_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_199_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10679_ _10679_/A vssd1 vssd1 vccd1 vccd1 _10679_/X sky130_fd_sc_hd__buf_2
X_15206_ _15239_/A _15206_/B vssd1 vssd1 vccd1 vccd1 _15206_/Y sky130_fd_sc_hd__nand2_1
XFILLER_199_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12418_ _12450_/B _12420_/C _17899_/Q vssd1 vssd1 vccd1 vccd1 _12419_/A sky130_fd_sc_hd__o21ai_2
X_16186_ _16188_/B _16183_/X _16184_/Y _16185_/X vssd1 vssd1 vccd1 vccd1 _18619_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_127_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13398_ _13398_/A vssd1 vssd1 vccd1 vccd1 _13398_/Y sky130_fd_sc_hd__inv_2
XFILLER_182_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_1295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15137_ _15142_/B _15135_/X _15136_/X _15123_/X vssd1 vssd1 vccd1 vccd1 _18372_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_127_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12349_ _17890_/Q _12340_/C _12184_/X vssd1 vssd1 vccd1 vccd1 _17890_/D sky130_fd_sc_hd__o21a_1
XFILLER_5_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15068_ _15247_/A vssd1 vssd1 vccd1 vccd1 _15115_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_4_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14019_ _14019_/A vssd1 vssd1 vccd1 vccd1 _14019_/X sky130_fd_sc_hd__buf_8
XFILLER_4_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_228_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_110_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_229_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18827_ _18860_/CLK _18827_/D vssd1 vssd1 vccd1 vccd1 _18827_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_3_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09560_ _09560_/A vssd1 vssd1 vccd1 vccd1 _09598_/S sky130_fd_sc_hd__buf_2
XFILLER_95_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18758_ _18786_/CLK _18758_/D vssd1 vssd1 vccd1 vccd1 _18758_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_209_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_1368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17709_ _17709_/A _17709_/B vssd1 vssd1 vccd1 vccd1 _17710_/A sky130_fd_sc_hd__or2_1
X_09491_ _18188_/Q _18187_/Q _18186_/Q _18185_/Q vssd1 vssd1 vccd1 vccd1 _13357_/B
+ sky130_fd_sc_hd__nor4_4
XFILLER_70_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18689_ _18693_/CLK _18689_/D vssd1 vssd1 vccd1 vccd1 _18689_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_91_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_224_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_169_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_191_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_136_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_219_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_219_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09827_ _17781_/Q vssd1 vssd1 vccd1 vccd1 _09828_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_115_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_231_wb_clk_i clkbuf_5_0_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17907_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_228_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_230_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09758_ _18107_/Q _10611_/B _09757_/X vssd1 vssd1 vccd1 vccd1 _09760_/B sky130_fd_sc_hd__a21oi_1
XFILLER_206_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_228_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09689_ _12059_/A vssd1 vssd1 vccd1 vccd1 _09689_/X sky130_fd_sc_hd__clkbuf_4
XTAP_2136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11720_ _11720_/A _11720_/B vssd1 vssd1 vccd1 vccd1 _11720_/Y sky130_fd_sc_hd__nor2_1
XFILLER_226_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11651_ _11651_/A _11651_/B vssd1 vssd1 vccd1 vccd1 _11651_/Y sky130_fd_sc_hd__nand2_1
XFILLER_70_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_230_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_1292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10602_ _10291_/X _10599_/X _10601_/X _09974_/A vssd1 vssd1 vccd1 vccd1 _10602_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_23_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14370_ _14375_/B vssd1 vssd1 vccd1 vccd1 _14370_/Y sky130_fd_sc_hd__inv_2
XFILLER_70_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11582_ _11582_/A _11786_/B vssd1 vssd1 vccd1 vccd1 _11795_/B sky130_fd_sc_hd__nand2_1
XFILLER_80_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_211_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_195_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13321_ _13313_/X _13319_/X _13320_/Y vssd1 vssd1 vccd1 vccd1 _18091_/D sky130_fd_sc_hd__a21oi_1
XFILLER_127_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10533_ _10547_/A _10533_/B vssd1 vssd1 vccd1 vccd1 _10533_/Y sky130_fd_sc_hd__nor2_1
XFILLER_167_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_202_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16040_ _16039_/B _16038_/X _16039_/Y _16028_/X vssd1 vssd1 vccd1 vccd1 _18587_/D
+ sky130_fd_sc_hd__o211a_1
X_13252_ _13252_/A vssd1 vssd1 vccd1 vccd1 _18079_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_196_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10464_ _10559_/S vssd1 vssd1 vccd1 vccd1 _10464_/X sky130_fd_sc_hd__buf_4
XFILLER_108_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12203_ _11704_/C _12200_/X _12202_/Y _11863_/X vssd1 vssd1 vccd1 vccd1 _17850_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_182_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_159_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13183_ _13183_/A vssd1 vssd1 vccd1 vccd1 _18048_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_123_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10395_ _10605_/B _10380_/X _10394_/X _09981_/A vssd1 vssd1 vccd1 vccd1 _10395_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_135_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12134_ _12106_/X _12107_/Y _12120_/Y _12132_/X _12133_/Y vssd1 vssd1 vccd1 vccd1
+ _12134_/X sky130_fd_sc_hd__a2111o_1
XFILLER_150_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17991_ _18151_/CLK _17991_/D vssd1 vssd1 vccd1 vccd1 _17991_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_97_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16942_ _18836_/Q _18800_/Q _16947_/S vssd1 vssd1 vccd1 vccd1 _16942_/X sky130_fd_sc_hd__mux2_1
X_12065_ _12065_/A _12129_/A vssd1 vssd1 vccd1 vccd1 _12067_/B sky130_fd_sc_hd__xor2_1
XFILLER_145_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_1271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11016_ _13375_/B _13375_/C _11037_/C vssd1 vssd1 vccd1 vccd1 _11017_/A sky130_fd_sc_hd__and3b_1
XFILLER_133_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16873_ _18821_/Q _18785_/Q _16900_/S vssd1 vssd1 vccd1 vccd1 _16873_/X sky130_fd_sc_hd__mux2_1
XFILLER_49_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18612_ _18614_/CLK _18612_/D vssd1 vssd1 vccd1 vccd1 _18612_/Q sky130_fd_sc_hd__dfxtp_2
X_15824_ _18534_/Q _15829_/B _15822_/X _15823_/X vssd1 vssd1 vccd1 vccd1 _18534_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_4050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_231_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_219_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_225_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18543_ _18582_/CLK _18543_/D vssd1 vssd1 vccd1 vccd1 _18543_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_4094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15755_ _15754_/B _15753_/X _15754_/Y _15740_/X vssd1 vssd1 vccd1 vccd1 _18518_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_3360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12967_ _12967_/A _12983_/A vssd1 vssd1 vccd1 vccd1 _12969_/C sky130_fd_sc_hd__xnor2_1
XFILLER_52_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14706_ _15145_/C _14706_/B vssd1 vssd1 vccd1 vccd1 _14772_/A sky130_fd_sc_hd__or2_1
XFILLER_61_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11918_ _11918_/A _11918_/B vssd1 vssd1 vccd1 vccd1 _11919_/B sky130_fd_sc_hd__xnor2_2
XFILLER_209_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18474_ _18506_/CLK _18474_/D vssd1 vssd1 vccd1 vccd1 _18474_/Q sky130_fd_sc_hd__dfxtp_1
X_15686_ _18537_/Q _18501_/Q _15693_/S vssd1 vssd1 vccd1 vccd1 _15686_/X sky130_fd_sc_hd__mux2_1
XFILLER_61_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12898_ _12898_/A vssd1 vssd1 vccd1 vccd1 _17962_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17425_ _17437_/A _17425_/B _17460_/C vssd1 vssd1 vccd1 vccd1 _17425_/X sky130_fd_sc_hd__or3_1
X_11849_ _11663_/X _11848_/X _11845_/A vssd1 vssd1 vccd1 vccd1 _11850_/D sky130_fd_sc_hd__a21oi_1
X_14637_ _14637_/A _14660_/B vssd1 vssd1 vccd1 vccd1 _16905_/A sky130_fd_sc_hd__or2_4
XFILLER_92_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_193_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14568_ _16835_/A vssd1 vssd1 vccd1 vccd1 _16839_/A sky130_fd_sc_hd__buf_8
XFILLER_18_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17356_ _18937_/Q _18901_/Q _17367_/S vssd1 vssd1 vccd1 vccd1 _17356_/X sky130_fd_sc_hd__mux2_1
XFILLER_105_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_220_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_35_wb_clk_i clkbuf_5_7_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18845_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_16307_ _16745_/A _16307_/B vssd1 vssd1 vccd1 vccd1 _16317_/B sky130_fd_sc_hd__nor2_1
XFILLER_53_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13519_ _13552_/B _13557_/A vssd1 vssd1 vccd1 vccd1 _13741_/A sky130_fd_sc_hd__nor2_1
XFILLER_119_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14499_ _14499_/A vssd1 vssd1 vccd1 vccd1 _18223_/D sky130_fd_sc_hd__clkbuf_1
X_17287_ _17334_/A _17291_/B vssd1 vssd1 vccd1 vccd1 _17287_/Y sky130_fd_sc_hd__nand2_1
XFILLER_220_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19026_ _19026_/CLK _19026_/D vssd1 vssd1 vccd1 vccd1 _19026_/Q sky130_fd_sc_hd__dfxtp_1
X_16238_ _16243_/B _16236_/X _16237_/X _16230_/X vssd1 vssd1 vccd1 vccd1 _18630_/D
+ sky130_fd_sc_hd__o211a_1
X_16169_ _16175_/B _16166_/X _16168_/X _16162_/X vssd1 vssd1 vccd1 vccd1 _18615_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_170_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08991_ _08991_/A vssd1 vssd1 vccd1 vccd1 _08991_/Y sky130_fd_sc_hd__inv_2
XFILLER_88_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_1322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_228_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09612_ _10110_/A vssd1 vssd1 vccd1 vccd1 _12056_/A sky130_fd_sc_hd__buf_2
XFILLER_216_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_228_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09543_ _18125_/Q _09530_/B _09530_/A vssd1 vssd1 vccd1 vccd1 _09560_/A sky130_fd_sc_hd__a21bo_2
XFILLER_83_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_221_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_221_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09474_ _09474_/A vssd1 vssd1 vccd1 vccd1 _09474_/Y sky130_fd_sc_hd__inv_2
XFILLER_212_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_212_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_197_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_184_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_212_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_211_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_137_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_180_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_133_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10180_ _10939_/B _12047_/A vssd1 vssd1 vccd1 vccd1 _10271_/B sky130_fd_sc_hd__and2_1
XFILLER_117_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_219_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13870_ _18460_/Q _13588_/A _13861_/A _18475_/Q vssd1 vssd1 vccd1 vccd1 _13870_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_101_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_219_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_207_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12821_ _12570_/B _12816_/X _12824_/A _12630_/B _12820_/X vssd1 vssd1 vccd1 vccd1
+ _12821_/Y sky130_fd_sc_hd__o221ai_1
XFILLER_76_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_215_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15540_ _15551_/A _15984_/B _15574_/C vssd1 vssd1 vccd1 vccd1 _15540_/X sky130_fd_sc_hd__or3_1
X_12752_ _12752_/A _12752_/B _12752_/C vssd1 vssd1 vccd1 vccd1 _12921_/B sky130_fd_sc_hd__and3_1
XTAP_1210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_1204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11703_ _11703_/A vssd1 vssd1 vccd1 vccd1 _11704_/B sky130_fd_sc_hd__inv_2
X_15471_ _15508_/A _15473_/B vssd1 vssd1 vccd1 vccd1 _15471_/Y sky130_fd_sc_hd__nand2_1
XTAP_1254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_203_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12683_ _12707_/A _17934_/Q vssd1 vssd1 vccd1 vccd1 _12688_/A sky130_fd_sc_hd__xnor2_1
XTAP_1276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_231_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_203_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14422_ _14422_/A vssd1 vssd1 vccd1 vccd1 _14422_/X sky130_fd_sc_hd__clkbuf_2
X_17210_ _17210_/A _17213_/B vssd1 vssd1 vccd1 vccd1 _17210_/Y sky130_fd_sc_hd__nand2_1
X_11634_ _11253_/A _11499_/B _11257_/B _11609_/A _11764_/A vssd1 vssd1 vccd1 vccd1
+ _11635_/C sky130_fd_sc_hd__o32a_1
X_18190_ _18960_/CLK _18190_/D vssd1 vssd1 vccd1 vccd1 _18190_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_156_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_196_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14353_ _17575_/A vssd1 vssd1 vccd1 vccd1 _14584_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_17141_ _17143_/B _17138_/X _17139_/Y _17140_/X vssd1 vssd1 vccd1 vccd1 _18847_/D
+ sky130_fd_sc_hd__o211a_1
X_11565_ _19032_/Q _11565_/B _12267_/A vssd1 vssd1 vccd1 vccd1 _11565_/X sky130_fd_sc_hd__and3_1
XFILLER_144_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13304_ _13304_/A _13304_/B vssd1 vssd1 vccd1 vccd1 _13311_/C sky130_fd_sc_hd__or2_1
XFILLER_6_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17072_ _17072_/A _17506_/B _17085_/C vssd1 vssd1 vccd1 vccd1 _17072_/X sky130_fd_sc_hd__or3_1
X_10516_ _10461_/X _10482_/X _10502_/X _10515_/X vssd1 vssd1 vccd1 vccd1 _10516_/Y
+ sky130_fd_sc_hd__a22oi_1
XFILLER_196_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14284_ _18175_/Q vssd1 vssd1 vccd1 vccd1 _15607_/B sky130_fd_sc_hd__buf_2
X_11496_ _11496_/A vssd1 vssd1 vccd1 vccd1 _11496_/Y sky130_fd_sc_hd__inv_2
XFILLER_6_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16023_ _18619_/Q _18583_/Q _16031_/S vssd1 vssd1 vccd1 vccd1 _16023_/X sky130_fd_sc_hd__mux2_1
X_13235_ _13257_/A vssd1 vssd1 vccd1 vccd1 _13244_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_108_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10447_ _10445_/X _10446_/X _10496_/A vssd1 vssd1 vccd1 vccd1 _10447_/X sky130_fd_sc_hd__mux2_1
XFILLER_109_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_226_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13166_ _13199_/A vssd1 vssd1 vccd1 vccd1 _13175_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_3_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10378_ _09959_/X _10375_/X _10377_/X _10333_/S vssd1 vssd1 vccd1 vccd1 _10378_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_48_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12117_ _12117_/A _12117_/B vssd1 vssd1 vccd1 vccd1 _12118_/B sky130_fd_sc_hd__xnor2_1
Xclkbuf_leaf_153_wb_clk_i _18102_/CLK vssd1 vssd1 vccd1 vccd1 _18110_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_112_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13097_ _16891_/A vssd1 vssd1 vccd1 vccd1 _13142_/A sky130_fd_sc_hd__clkbuf_2
X_17974_ _19027_/CLK _17974_/D vssd1 vssd1 vccd1 vccd1 _17974_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_97_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16925_ _18832_/Q _18796_/Q _16925_/S vssd1 vssd1 vccd1 vccd1 _16925_/X sky130_fd_sc_hd__mux2_1
X_12048_ _12048_/A vssd1 vssd1 vccd1 vccd1 _12055_/A sky130_fd_sc_hd__buf_4
XFILLER_172_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16856_ _18817_/Q _18781_/Q _16864_/S vssd1 vssd1 vccd1 vccd1 _16856_/X sky130_fd_sc_hd__mux2_1
XFILLER_20_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15807_ _15806_/B _15805_/X _15806_/Y _15803_/X vssd1 vssd1 vccd1 vccd1 _18530_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_225_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16787_ _16787_/A vssd1 vssd1 vccd1 vccd1 _16802_/S sky130_fd_sc_hd__clkbuf_2
X_13999_ _18589_/Q _13730_/A _13780_/A _18580_/Q _13998_/X vssd1 vssd1 vccd1 vccd1
+ _13999_/X sky130_fd_sc_hd__a221o_1
XFILLER_46_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18526_ _18563_/CLK _18526_/D vssd1 vssd1 vccd1 vccd1 _18526_/Q sky130_fd_sc_hd__dfxtp_4
X_15738_ _15751_/A _15743_/B vssd1 vssd1 vccd1 vccd1 _15738_/Y sky130_fd_sc_hd__nand2_1
XFILLER_94_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_222_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_222_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_1318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18457_ _18458_/CLK _18457_/D vssd1 vssd1 vccd1 vccd1 _18457_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_178_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15669_ _18532_/Q _18496_/Q _15693_/S vssd1 vssd1 vccd1 vccd1 _15669_/X sky130_fd_sc_hd__mux2_1
XFILLER_205_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17408_ _17456_/A _17408_/B vssd1 vssd1 vccd1 vccd1 _17408_/Y sky130_fd_sc_hd__nand2_1
X_09190_ _18581_/Q _18580_/Q _18579_/Q vssd1 vssd1 vccd1 vccd1 _09193_/B sky130_fd_sc_hd__or3_4
XFILLER_92_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18388_ _18398_/CLK _18388_/D vssd1 vssd1 vccd1 vccd1 _18388_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_21_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_187_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17339_ _18933_/Q _18897_/Q _17347_/S vssd1 vssd1 vccd1 vccd1 _17339_/X sky130_fd_sc_hd__mux2_1
XFILLER_174_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_119_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_220_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19009_ _19009_/CLK _19009_/D vssd1 vssd1 vccd1 vccd1 _19009_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_161_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_216_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08974_ _08998_/A vssd1 vssd1 vccd1 vccd1 _08979_/A sky130_fd_sc_hd__buf_12
XTAP_5509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_1283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_227_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09526_ _14299_/A vssd1 vssd1 vccd1 vccd1 _14222_/A sky130_fd_sc_hd__buf_4
XFILLER_71_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_212_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_197_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_227_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_213_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_212_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09457_ _18134_/D _09457_/B vssd1 vssd1 vccd1 vccd1 _09458_/A sky130_fd_sc_hd__or2_4
XPHY_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_227_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09388_ _18371_/Q _18370_/Q _18369_/Q vssd1 vssd1 vccd1 vccd1 _09952_/A sky130_fd_sc_hd__or3_4
XFILLER_138_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_196_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_177_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11350_ _11442_/A _11455_/C vssd1 vssd1 vccd1 vccd1 _11495_/D sky130_fd_sc_hd__and2b_1
XFILLER_180_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_117_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10301_ _10278_/A _10299_/X _10300_/X _09976_/A vssd1 vssd1 vccd1 vccd1 _10301_/X
+ sky130_fd_sc_hd__a22o_1
X_11281_ _11281_/A _11281_/B _13443_/A _11280_/Y vssd1 vssd1 vccd1 vccd1 _11281_/X
+ sky130_fd_sc_hd__or4b_1
XFILLER_106_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13020_ _13039_/B vssd1 vssd1 vccd1 vccd1 _13036_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_193_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10232_ _10232_/A _10232_/B vssd1 vssd1 vccd1 vccd1 _10521_/A sky130_fd_sc_hd__xnor2_4
XFILLER_134_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_180_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_121_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10163_ _10133_/A _10175_/A _10178_/A _10178_/B vssd1 vssd1 vccd1 vccd1 _10172_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_79_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14971_ _14995_/A _14971_/B vssd1 vssd1 vccd1 vccd1 _14971_/Y sky130_fd_sc_hd__nand2_1
X_10094_ _09277_/A _09277_/B _09277_/C _09277_/D _10955_/S _09987_/X vssd1 vssd1 vccd1
+ vccd1 _10094_/X sky130_fd_sc_hd__mux4_1
XFILLER_130_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16710_ _18782_/Q _18746_/Q _16715_/S vssd1 vssd1 vccd1 vccd1 _16710_/X sky130_fd_sc_hd__mux2_1
XFILLER_48_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13922_ _18742_/Q _13619_/A _13918_/X _13921_/X vssd1 vssd1 vccd1 vccd1 _13922_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_43_1277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17690_ _17712_/A _17690_/B vssd1 vssd1 vccd1 vccd1 _17691_/A sky130_fd_sc_hd__and2_1
XFILLER_101_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16641_ _16641_/A vssd1 vssd1 vccd1 vccd1 _16657_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_63_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13853_ _18730_/Q _13551_/X _13851_/X _13852_/X vssd1 vssd1 vccd1 vccd1 _13853_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_142_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12804_ _12699_/Y _17967_/Q _12542_/B _12846_/A vssd1 vssd1 vccd1 vccd1 _12804_/X
+ sky130_fd_sc_hd__o2bb2a_1
X_16572_ _16572_/A _16575_/B vssd1 vssd1 vccd1 vccd1 _16572_/Y sky130_fd_sc_hd__nand2_1
XFILLER_16_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_188_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13784_ _18414_/Q _13642_/A _13764_/X _18438_/Q vssd1 vssd1 vccd1 vccd1 _13784_/X
+ sky130_fd_sc_hd__a22o_1
X_10996_ _18994_/Q _10977_/X _10990_/X vssd1 vssd1 vccd1 vccd1 _18994_/D sky130_fd_sc_hd__a21bo_1
XFILLER_204_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_215_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18311_ _18312_/CLK _18311_/D vssd1 vssd1 vccd1 vccd1 _18311_/Q sky130_fd_sc_hd__dfxtp_4
X_15523_ _18497_/Q _18461_/Q _15545_/S vssd1 vssd1 vccd1 vccd1 _15523_/X sky130_fd_sc_hd__mux2_1
XTAP_1040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_187_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12735_ _19016_/Q _19015_/Q _19018_/Q _19017_/Q vssd1 vssd1 vccd1 vccd1 _12736_/C
+ sky130_fd_sc_hd__and4_1
XFILLER_35_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_203_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_206_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_230_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_231_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18242_ _18245_/CLK _18242_/D vssd1 vssd1 vccd1 vccd1 _18242_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15454_ _18481_/Q _18445_/Q _15458_/S vssd1 vssd1 vccd1 vccd1 _15454_/X sky130_fd_sc_hd__mux2_1
XTAP_1095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12666_ _12665_/A _12665_/B _12591_/X vssd1 vssd1 vccd1 vccd1 _12666_/X sky130_fd_sc_hd__o21a_1
XFILLER_31_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11617_ _11617_/A _11617_/B _11617_/C _11546_/A vssd1 vssd1 vccd1 vccd1 _11617_/X
+ sky130_fd_sc_hd__or4b_2
X_14405_ _14423_/A vssd1 vssd1 vccd1 vccd1 _14405_/X sky130_fd_sc_hd__clkbuf_2
X_18173_ _18178_/CLK _18173_/D vssd1 vssd1 vccd1 vccd1 _18173_/Q sky130_fd_sc_hd__dfxtp_1
X_15385_ _15578_/A vssd1 vssd1 vccd1 vccd1 _15442_/A sky130_fd_sc_hd__clkbuf_2
X_12597_ _17927_/Q _12597_/B vssd1 vssd1 vccd1 vccd1 _12598_/B sky130_fd_sc_hd__nor2_1
XFILLER_15_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17124_ _17254_/B vssd1 vssd1 vccd1 vccd1 _17173_/C sky130_fd_sc_hd__clkbuf_2
X_11548_ _11495_/B _11354_/B _11547_/Y _11683_/A vssd1 vssd1 vccd1 vccd1 _11844_/A
+ sky130_fd_sc_hd__o211a_1
X_14336_ _14325_/A _14335_/X _14222_/A vssd1 vssd1 vccd1 vccd1 _14336_/X sky130_fd_sc_hd__a21o_1
XFILLER_128_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_143_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17055_ _18863_/Q _18827_/Q _17055_/S vssd1 vssd1 vccd1 vccd1 _17055_/X sky130_fd_sc_hd__mux2_1
XFILLER_13_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14267_ _14267_/A _14267_/B vssd1 vssd1 vccd1 vccd1 _14267_/Y sky130_fd_sc_hd__nand2_1
X_11479_ _17887_/Q _11479_/B vssd1 vssd1 vccd1 vccd1 _11489_/B sky130_fd_sc_hd__or2_1
XFILLER_125_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16006_ _18615_/Q _18579_/Q _16010_/S vssd1 vssd1 vccd1 vccd1 _16006_/X sky130_fd_sc_hd__mux2_1
X_13218_ _13222_/A _18065_/Q vssd1 vssd1 vccd1 vccd1 _13219_/A sky130_fd_sc_hd__and2_1
XFILLER_131_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14198_ _18211_/Q _14470_/A _14192_/X _14216_/B _14216_/A vssd1 vssd1 vccd1 vccd1
+ _14349_/B sky130_fd_sc_hd__a311o_2
XFILLER_98_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_112_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13149_ _13151_/A _18034_/Q vssd1 vssd1 vccd1 vccd1 _13150_/A sky130_fd_sc_hd__and2_1
XTAP_835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17957_ _17959_/CLK _17957_/D vssd1 vssd1 vccd1 vccd1 _17957_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_97_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_1366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16908_ _18828_/Q _18792_/Q _16925_/S vssd1 vssd1 vccd1 vccd1 _16908_/X sky130_fd_sc_hd__mux2_1
XFILLER_78_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17888_ _17888_/CLK _17888_/D vssd1 vssd1 vccd1 vccd1 _17888_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_26_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16839_ _16839_/A vssd1 vssd1 vccd1 vccd1 _17437_/B sky130_fd_sc_hd__buf_4
XFILLER_38_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_202_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_50_wb_clk_i clkbuf_5_16_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18826_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_09311_ _18479_/Q _18478_/Q _18477_/Q vssd1 vssd1 vccd1 vccd1 _09314_/B sky130_fd_sc_hd__or3_2
XFILLER_34_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_222_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_206_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18509_ _18546_/CLK _18509_/D vssd1 vssd1 vccd1 vccd1 _18509_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_202_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_178_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09242_ _18914_/Q _18913_/Q _18912_/Q vssd1 vssd1 vccd1 vccd1 _09243_/D sky130_fd_sc_hd__or3_4
XFILLER_221_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09173_ _18626_/Q _18625_/Q _18624_/Q vssd1 vssd1 vccd1 vccd1 _09176_/B sky130_fd_sc_hd__or3_4
XFILLER_181_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_222_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_192_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08957_ _08960_/A vssd1 vssd1 vccd1 vccd1 _08957_/Y sky130_fd_sc_hd__inv_2
XTAP_4605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10850_ _10616_/Y _10709_/X _10752_/X _10849_/X vssd1 vssd1 vccd1 vccd1 _10850_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_60_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09509_ _12972_/A _09518_/B vssd1 vssd1 vccd1 vccd1 _09509_/Y sky130_fd_sc_hd__nor2_2
XPHY_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10781_ _09332_/A _09337_/B _10781_/S vssd1 vssd1 vccd1 vccd1 _10781_/X sky130_fd_sc_hd__mux2_1
XFILLER_25_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_112_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_212_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12520_ _13153_/A _12520_/B vssd1 vssd1 vccd1 vccd1 _17915_/D sky130_fd_sc_hd__nor2_1
XFILLER_200_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_201_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12451_ _12458_/A _12451_/B vssd1 vssd1 vccd1 vccd1 _12452_/C sky130_fd_sc_hd__nand2_1
X_11402_ _17796_/Q _17797_/Q _17798_/Q vssd1 vssd1 vccd1 vccd1 _11497_/B sky130_fd_sc_hd__o21a_2
X_15170_ _15169_/B _15168_/X _15169_/Y _15166_/X vssd1 vssd1 vccd1 vccd1 _18380_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_138_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12382_ _12373_/A _18987_/Q _18105_/Q vssd1 vssd1 vccd1 vccd1 _12384_/C sky130_fd_sc_hd__o21a_1
XFILLER_197_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14121_ _18902_/Q _13562_/A _13858_/X _18893_/Q vssd1 vssd1 vccd1 vccd1 _14121_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_158_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11333_ _11333_/A vssd1 vssd1 vccd1 vccd1 _11333_/Y sky130_fd_sc_hd__inv_2
XFILLER_125_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14052_ _18500_/Q _13877_/X _13842_/A _18494_/Q _14051_/X vssd1 vssd1 vccd1 vccd1
+ _14052_/X sky130_fd_sc_hd__a221o_1
XFILLER_4_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11264_ _12037_/A vssd1 vssd1 vccd1 vccd1 _11264_/Y sky130_fd_sc_hd__inv_2
XFILLER_98_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_1344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13003_ _13000_/A _12991_/X _13002_/X _12964_/X vssd1 vssd1 vccd1 vccd1 _17980_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_180_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10215_ _10215_/A _10215_/B vssd1 vssd1 vccd1 vccd1 _10227_/B sky130_fd_sc_hd__xnor2_4
Xclkbuf_2_3_0_wb_clk_i clkbuf_2_3_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_2_3_1_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_140_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18860_ _18860_/CLK _18860_/D vssd1 vssd1 vccd1 vccd1 _18860_/Q sky130_fd_sc_hd__dfxtp_2
X_11195_ _11195_/A vssd1 vssd1 vccd1 vccd1 _17810_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_79_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17811_ _17851_/CLK _17811_/D vssd1 vssd1 vccd1 vccd1 _17811_/Q sky130_fd_sc_hd__dfxtp_1
X_10146_ _10146_/A _10146_/B vssd1 vssd1 vccd1 vccd1 _10147_/B sky130_fd_sc_hd__and2_1
X_18791_ _18823_/CLK _18791_/D vssd1 vssd1 vccd1 vccd1 _18791_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_94_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17742_ _17742_/A vssd1 vssd1 vccd1 vccd1 _19014_/D sky130_fd_sc_hd__clkbuf_1
XTAP_5873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14954_ _14960_/B _14952_/X _14953_/X _14941_/X vssd1 vssd1 vccd1 vccd1 _18327_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_48_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10077_ _10966_/B _10073_/X _10076_/X _09728_/D vssd1 vssd1 vccd1 vccd1 _10077_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_5884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_1366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13905_ _13899_/X _13901_/X _13904_/X _13684_/Y vssd1 vssd1 vccd1 vccd1 _13905_/X
+ sky130_fd_sc_hd__o31a_1
XFILLER_208_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17673_ _17673_/A vssd1 vssd1 vccd1 vccd1 _18980_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_208_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14885_ _14932_/A _14890_/B vssd1 vssd1 vccd1 vccd1 _14885_/Y sky130_fd_sc_hd__nand2_1
XFILLER_223_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16624_ _16623_/B _16622_/X _16623_/Y _16619_/X vssd1 vssd1 vccd1 vccd1 _18725_/D
+ sky130_fd_sc_hd__o211a_1
XINSDIODE2_203 _12346_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13836_ _18685_/Q _13621_/X _13834_/X _18679_/Q _13835_/X vssd1 vssd1 vccd1 vccd1
+ _13836_/X sky130_fd_sc_hd__a221o_1
XINSDIODE2_214 _13654_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_169_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XINSDIODE2_225 _15643_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XINSDIODE2_236 input1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_247 _08954_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16555_ _16555_/A _16703_/B _16568_/C vssd1 vssd1 vccd1 vccd1 _16555_/X sky130_fd_sc_hd__or3_1
XINSDIODE2_258 _13612_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13767_ _18501_/Q _13742_/X _13766_/X _18483_/Q vssd1 vssd1 vccd1 vccd1 _13767_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_44_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10979_ input2/X vssd1 vssd1 vccd1 vccd1 _12361_/A sky130_fd_sc_hd__buf_6
XFILLER_62_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_269 _18425_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15506_ _15511_/B _15503_/X _15505_/X _15496_/X vssd1 vssd1 vccd1 vccd1 _18456_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_31_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12718_ _12962_/A vssd1 vssd1 vccd1 vccd1 _12718_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_188_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16486_ _18728_/Q _18692_/Q _16490_/S vssd1 vssd1 vccd1 vccd1 _16486_/X sky130_fd_sc_hd__mux2_1
XFILLER_31_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13698_ _13698_/A vssd1 vssd1 vccd1 vccd1 _14026_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_30_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18225_ _19026_/CLK _18225_/D vssd1 vssd1 vccd1 vccd1 _18225_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15437_ _16949_/A vssd1 vssd1 vccd1 vccd1 _16032_/B sky130_fd_sc_hd__buf_2
XFILLER_175_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12649_ _12649_/A _12649_/B vssd1 vssd1 vccd1 vccd1 _12649_/Y sky130_fd_sc_hd__nand2_1
XFILLER_191_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18156_ _18163_/CLK _18156_/D vssd1 vssd1 vccd1 vccd1 _18156_/Q sky130_fd_sc_hd__dfxtp_1
X_15368_ _15527_/A _15451_/C vssd1 vssd1 vccd1 vccd1 _15375_/B sky130_fd_sc_hd__nor2_1
XFILLER_191_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17107_ _17536_/A _17107_/B vssd1 vssd1 vccd1 vccd1 _17115_/B sky130_fd_sc_hd__nor2_1
XFILLER_190_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14319_ _14318_/X _12133_/A _14319_/S vssd1 vssd1 vccd1 vccd1 _14321_/B sky130_fd_sc_hd__mux2_1
XFILLER_171_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18087_ _18087_/CLK _18087_/D vssd1 vssd1 vccd1 vccd1 _18087_/Q sky130_fd_sc_hd__dfxtp_1
X_15299_ _15358_/A _15909_/B _15358_/C vssd1 vssd1 vccd1 vccd1 _15299_/X sky130_fd_sc_hd__or3_1
X_19125__96 vssd1 vssd1 vccd1 vccd1 _19125__96/HI _19233_/A sky130_fd_sc_hd__conb_1
XFILLER_7_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17038_ _17107_/B vssd1 vssd1 vccd1 vccd1 _17085_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_104_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_217_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09860_ _09860_/A _09860_/B _09860_/C vssd1 vssd1 vccd1 vccd1 _09862_/A sky130_fd_sc_hd__nor3_2
XFILLER_124_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09791_ _09892_/A _09789_/X _09790_/X vssd1 vssd1 vccd1 vccd1 _09813_/A sky130_fd_sc_hd__a21o_1
XTAP_665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18989_ _18989_/CLK _18989_/D vssd1 vssd1 vccd1 vccd1 _18989_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_85_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_227_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_227_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_1366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_226_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_1264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_1215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_226_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_214_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_1305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_224_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09225_ _18938_/Q _18937_/Q _18936_/Q vssd1 vssd1 vccd1 vccd1 _09227_/C sky130_fd_sc_hd__or3_2
XFILLER_158_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_210_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09156_ _18653_/Q _18652_/Q _18651_/Q vssd1 vssd1 vccd1 vccd1 _09160_/A sky130_fd_sc_hd__or3_4
XFILLER_154_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09087_ _17838_/Q _17837_/Q _17836_/Q vssd1 vssd1 vccd1 vccd1 _09088_/A sky130_fd_sc_hd__and3_1
XFILLER_68_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10000_ _10086_/A vssd1 vssd1 vccd1 vccd1 _10940_/A sky130_fd_sc_hd__buf_4
XFILLER_192_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09989_ _09148_/A _09143_/D _12059_/A vssd1 vssd1 vccd1 vccd1 _09989_/X sky130_fd_sc_hd__mux2_1
XTAP_5147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_218_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_229_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11951_ _11951_/A _11951_/B vssd1 vssd1 vccd1 vccd1 _11985_/A sky130_fd_sc_hd__xnor2_4
XFILLER_218_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_205_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10902_ _10900_/X _10901_/X _10902_/S vssd1 vssd1 vccd1 vccd1 _10902_/X sky130_fd_sc_hd__mux2_1
XFILLER_205_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14670_ _14683_/A _14670_/B vssd1 vssd1 vccd1 vccd1 _14670_/Y sky130_fd_sc_hd__nand2_1
XTAP_3778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11882_ hold4/X _11867_/X _11870_/Y vssd1 vssd1 vccd1 vccd1 _11883_/B sky130_fd_sc_hd__a21oi_1
XTAP_3789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_189_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13621_ _13621_/A vssd1 vssd1 vccd1 vccd1 _13621_/X sky130_fd_sc_hd__buf_6
XFILLER_72_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10833_ _10833_/A _10833_/B _10833_/C vssd1 vssd1 vccd1 vccd1 _10833_/X sky130_fd_sc_hd__and3_1
XFILLER_32_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_198_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16340_ _18692_/Q _18656_/Q _16345_/S vssd1 vssd1 vccd1 vccd1 _16340_/X sky130_fd_sc_hd__mux2_1
X_13552_ _13563_/A _13552_/B vssd1 vssd1 vccd1 vccd1 _13906_/B sky130_fd_sc_hd__nor2_4
X_10764_ _10764_/A _10764_/B vssd1 vssd1 vccd1 vccd1 _10764_/X sky130_fd_sc_hd__or2_1
XFILLER_164_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12503_ _17911_/Q _12501_/X _12502_/Y vssd1 vssd1 vccd1 vccd1 _17911_/D sky130_fd_sc_hd__a21oi_1
XFILLER_12_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16271_ _18675_/Q _18639_/Q _16271_/S vssd1 vssd1 vccd1 vccd1 _16271_/X sky130_fd_sc_hd__mux2_1
XFILLER_186_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13483_ _14420_/A _13483_/B vssd1 vssd1 vccd1 vccd1 _18164_/D sky130_fd_sc_hd__nor2_1
X_10695_ _10695_/A vssd1 vssd1 vccd1 vccd1 _10695_/X sky130_fd_sc_hd__buf_4
X_18010_ _19004_/CLK _18010_/D vssd1 vssd1 vccd1 vccd1 _18010_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15222_ _18430_/Q _18394_/Q _15226_/S vssd1 vssd1 vccd1 vccd1 _15222_/X sky130_fd_sc_hd__mux2_1
XFILLER_12_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12434_ _12412_/A _12413_/X _12419_/A _12420_/X _12429_/A vssd1 vssd1 vccd1 vccd1
+ _12439_/D sky130_fd_sc_hd__o2111ai_2
XFILLER_201_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15153_ _18376_/Q _15154_/B _15152_/Y _15143_/X vssd1 vssd1 vccd1 vccd1 _18376_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_172_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12365_ _12373_/A _17893_/Q vssd1 vssd1 vccd1 vccd1 _12365_/X sky130_fd_sc_hd__or2b_2
XFILLER_148_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14104_ _18794_/Q _13848_/X _13702_/A _18788_/Q vssd1 vssd1 vccd1 vccd1 _14104_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_153_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11316_ _11375_/B _11316_/B vssd1 vssd1 vccd1 vccd1 _11340_/B sky130_fd_sc_hd__nor2_2
XFILLER_181_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15084_ _15082_/B _15081_/X _15082_/Y _15083_/X vssd1 vssd1 vccd1 vccd1 _18359_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_154_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12296_ _17874_/Q _13066_/B _12304_/A vssd1 vssd1 vccd1 vccd1 _12297_/A sky130_fd_sc_hd__and3_1
XFILLER_113_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14035_ _18266_/Q _13612_/X _14027_/X _18257_/Q _14034_/X vssd1 vssd1 vccd1 vccd1
+ _14035_/X sky130_fd_sc_hd__a221o_1
X_18912_ _18914_/CLK _18912_/D vssd1 vssd1 vccd1 vccd1 _18912_/Q sky130_fd_sc_hd__dfxtp_1
X_11247_ _11498_/A vssd1 vssd1 vccd1 vccd1 _13501_/A sky130_fd_sc_hd__inv_2
XFILLER_84_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18843_ _18845_/CLK _18843_/D vssd1 vssd1 vccd1 vccd1 _18843_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_68_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11178_ _11184_/C _11198_/B _11178_/C vssd1 vssd1 vccd1 vccd1 _11179_/A sky130_fd_sc_hd__and3b_1
XFILLER_79_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10129_ _10159_/A _10129_/B vssd1 vssd1 vccd1 vccd1 _10440_/B sky130_fd_sc_hd__xnor2_4
XFILLER_110_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18774_ _18799_/CLK _18774_/D vssd1 vssd1 vccd1 vccd1 _18774_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_83_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15986_ _18610_/Q _18574_/Q _15990_/S vssd1 vssd1 vccd1 vccd1 _15986_/X sky130_fd_sc_hd__mux2_1
XFILLER_48_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17725_ _17736_/A vssd1 vssd1 vccd1 vccd1 _17734_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_212_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14937_ _15229_/A _14937_/B vssd1 vssd1 vccd1 vccd1 _14949_/B sky130_fd_sc_hd__nor2_1
XFILLER_36_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17656_ _17659_/A _17656_/B vssd1 vssd1 vccd1 vccd1 _17657_/A sky130_fd_sc_hd__and2_1
X_14868_ _14928_/A vssd1 vssd1 vccd1 vccd1 _14919_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_1_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_224_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_223_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_224_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16607_ _18757_/Q _18721_/Q _16617_/S vssd1 vssd1 vccd1 vccd1 _16607_/X sky130_fd_sc_hd__mux2_1
X_13819_ _18945_/Q _13616_/A _13759_/A _18948_/Q _13818_/X vssd1 vssd1 vccd1 vccd1
+ _13819_/X sky130_fd_sc_hd__a221o_4
XFILLER_23_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17587_ _17587_/A _17587_/B vssd1 vssd1 vccd1 vccd1 _17588_/A sky130_fd_sc_hd__and2_1
X_14799_ _14881_/A vssd1 vssd1 vccd1 vccd1 _14799_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_91_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16538_ _16575_/A _16538_/B vssd1 vssd1 vccd1 vccd1 _16538_/Y sky130_fd_sc_hd__nand2_1
XFILLER_143_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16469_ _16475_/B _16467_/X _16468_/X _16456_/X vssd1 vssd1 vccd1 vccd1 _18687_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_177_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09010_ _09010_/A vssd1 vssd1 vccd1 vccd1 _09010_/Y sky130_fd_sc_hd__inv_2
X_18208_ _18992_/CLK _18208_/D vssd1 vssd1 vccd1 vccd1 _18208_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_223_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19188_ _19188_/A _09006_/Y vssd1 vssd1 vccd1 vccd1 io_out[26] sky130_fd_sc_hd__ebufn_8
XFILLER_191_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18139_ _18147_/CLK _18139_/D vssd1 vssd1 vccd1 vccd1 _18139_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_8_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09912_ _09953_/A vssd1 vssd1 vccd1 vccd1 _09959_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_137_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09843_ _09843_/A _09843_/B vssd1 vssd1 vccd1 vccd1 _09860_/A sky130_fd_sc_hd__xnor2_1
XFILLER_59_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09774_ _09774_/A _09774_/B vssd1 vssd1 vccd1 vccd1 _09918_/B sky130_fd_sc_hd__xnor2_4
XFILLER_26_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_230_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_214_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_199_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09208_ _18665_/Q _18664_/Q _18663_/Q vssd1 vssd1 vccd1 vccd1 _10795_/A sky130_fd_sc_hd__or3_4
XFILLER_139_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10480_ _10478_/X _10479_/X _10902_/S vssd1 vssd1 vccd1 vccd1 _10480_/X sky130_fd_sc_hd__mux2_1
XFILLER_136_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_202_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09139_ _18731_/Q _18730_/Q _18729_/Q vssd1 vssd1 vccd1 vccd1 _09993_/A sky130_fd_sc_hd__or3_4
XFILLER_154_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12150_ _12145_/A _12139_/A _12151_/A vssd1 vssd1 vccd1 vccd1 _12154_/B sky130_fd_sc_hd__mux2_1
XFILLER_162_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11101_ _11586_/A _17805_/Q _11113_/S vssd1 vssd1 vccd1 vccd1 _11102_/A sky130_fd_sc_hd__mux2_1
XFILLER_151_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12081_ _09684_/A _12079_/Y _12080_/X vssd1 vssd1 vccd1 vccd1 _12082_/B sky130_fd_sc_hd__o21ba_1
XFILLER_194_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11032_ _11032_/A _11031_/X vssd1 vssd1 vccd1 vccd1 _11038_/A sky130_fd_sc_hd__or2b_1
XFILLER_110_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_231_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_89_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_231_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15840_ _15840_/A vssd1 vssd1 vccd1 vccd1 _16273_/A sky130_fd_sc_hd__buf_2
XTAP_4210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15771_ _15915_/A _15894_/C vssd1 vssd1 vccd1 vccd1 _15782_/B sky130_fd_sc_hd__nor2_1
XTAP_4265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12983_ _12983_/A _12983_/B vssd1 vssd1 vccd1 vccd1 _12983_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_58_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17510_ _17512_/B _17508_/X _17509_/Y _17497_/X vssd1 vssd1 vccd1 vccd1 _18940_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_91_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14722_ _18306_/Q _18270_/Q _14736_/S vssd1 vssd1 vccd1 vccd1 _14722_/X sky130_fd_sc_hd__mux2_1
XTAP_3553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18490_ _18497_/CLK _18490_/D vssd1 vssd1 vccd1 vccd1 _18490_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_166_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11934_ _11963_/A vssd1 vssd1 vccd1 vccd1 _11934_/Y sky130_fd_sc_hd__clkinv_2
XTAP_3575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_178_wb_clk_i clkbuf_5_10_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18095_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_72_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17441_ _17497_/A vssd1 vssd1 vccd1 vccd1 _17441_/X sky130_fd_sc_hd__clkbuf_2
X_14653_ _16922_/A vssd1 vssd1 vccd1 vccd1 _15243_/B sky130_fd_sc_hd__buf_6
XFILLER_150_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11865_ _12224_/A vssd1 vssd1 vccd1 vccd1 _14421_/A sky130_fd_sc_hd__buf_4
XTAP_2874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_107_wb_clk_i clkbuf_5_29_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18572_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_13604_ _18828_/Q _13586_/A _13588_/A _18819_/Q vssd1 vssd1 vccd1 vccd1 _13604_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_60_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17372_ _17395_/A _17372_/B vssd1 vssd1 vccd1 vccd1 _17372_/Y sky130_fd_sc_hd__nand2_1
X_10816_ _10779_/X _10809_/X _10811_/X _10815_/X _10671_/B vssd1 vssd1 vccd1 vccd1
+ _10819_/B sky130_fd_sc_hd__a32o_1
X_14584_ _14584_/A _14584_/B _15186_/B vssd1 vssd1 vccd1 vccd1 _14584_/X sky130_fd_sc_hd__or3_1
XFILLER_14_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11796_ _11797_/A _11797_/B _11787_/X _11729_/X vssd1 vssd1 vccd1 vccd1 _11796_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_159_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_201_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16323_ _16329_/B _16320_/X _16322_/X _16314_/X vssd1 vssd1 vccd1 vccd1 _18651_/D
+ sky130_fd_sc_hd__o211a_1
X_13535_ _13535_/A vssd1 vssd1 vccd1 vccd1 _13706_/A sky130_fd_sc_hd__buf_4
XFILLER_41_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_207_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_203_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10747_ _10809_/A _10747_/B vssd1 vssd1 vccd1 vccd1 _10747_/X sky130_fd_sc_hd__or2_1
XFILLER_43_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16254_ _16327_/A vssd1 vssd1 vccd1 vccd1 _16271_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_9_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_186_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13466_ _17841_/Q _13464_/X _13465_/X vssd1 vssd1 vccd1 vccd1 _13467_/B sky130_fd_sc_hd__a21oi_1
X_10678_ _10867_/A vssd1 vssd1 vccd1 vccd1 _10678_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_199_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15205_ _18425_/Q _18389_/Q _15226_/S vssd1 vssd1 vccd1 vccd1 _15205_/X sky130_fd_sc_hd__mux2_1
XFILLER_138_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12417_ _18991_/Q _12426_/C vssd1 vssd1 vccd1 vccd1 _12420_/C sky130_fd_sc_hd__and2_1
X_16185_ _16252_/A vssd1 vssd1 vccd1 vccd1 _16185_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_154_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13397_ _18124_/Q _13336_/X _13395_/X vssd1 vssd1 vccd1 vccd1 _18124_/D sky130_fd_sc_hd__o21a_1
XFILLER_142_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_160_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15136_ _15162_/A _15279_/B _15136_/C vssd1 vssd1 vccd1 vccd1 _15136_/X sky130_fd_sc_hd__or3_1
XFILLER_142_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12348_ _12348_/A vssd1 vssd1 vccd1 vccd1 _17889_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_114_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15067_ _18354_/Q _15072_/B _15065_/X _15066_/X vssd1 vssd1 vccd1 vccd1 _18354_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_141_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12279_ _12279_/A _12279_/B vssd1 vssd1 vccd1 vccd1 _12279_/Y sky130_fd_sc_hd__nor2_1
XFILLER_4_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_214_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14018_ _18875_/Q _13838_/X _14017_/X _18851_/Q vssd1 vssd1 vccd1 vccd1 _14018_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_68_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_136_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_228_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18826_ _18826_/CLK _18826_/D vssd1 vssd1 vccd1 vccd1 _18826_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_56_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_110_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_209_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18757_ _18786_/CLK _18757_/D vssd1 vssd1 vccd1 vccd1 _18757_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_110_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15969_ _15971_/B _15967_/X _15968_/Y _15948_/X vssd1 vssd1 vccd1 vccd1 _18568_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_49_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17708_ _17779_/Q _09509_/Y _13363_/Y _18991_/Q vssd1 vssd1 vccd1 vccd1 _18991_/D
+ sky130_fd_sc_hd__a22o_1
X_09490_ _13416_/A vssd1 vssd1 vccd1 vccd1 _14297_/A sky130_fd_sc_hd__buf_4
X_18688_ _18693_/CLK _18688_/D vssd1 vssd1 vccd1 vccd1 _18688_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_110_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17639_ _17639_/A vssd1 vssd1 vccd1 vccd1 _18972_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_212_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_224_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_225_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_191_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_145_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_219_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09826_ _17975_/Q _17781_/Q vssd1 vssd1 vccd1 vccd1 _09834_/B sky130_fd_sc_hd__xor2_4
XFILLER_47_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_219_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09757_ _18096_/Q _13000_/C vssd1 vssd1 vccd1 vccd1 _09757_/X sky130_fd_sc_hd__and2_1
Xclkbuf_leaf_5_wb_clk_i _17929_/CLK vssd1 vssd1 vccd1 vccd1 _18196_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_230_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_230_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09688_ _09688_/A vssd1 vssd1 vccd1 vccd1 _12059_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_55_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_214_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_214_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_199_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11650_ _11642_/X _11645_/X _12253_/A _11649_/X _11689_/A vssd1 vssd1 vccd1 vccd1
+ _11651_/B sky130_fd_sc_hd__a32o_1
XTAP_1458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_230_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_211_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10601_ _09958_/A _09677_/X _10600_/X _10294_/X vssd1 vssd1 vccd1 vccd1 _10601_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_120_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11581_ _11617_/A _11788_/B vssd1 vssd1 vccd1 vccd1 _11786_/B sky130_fd_sc_hd__or2_1
XFILLER_195_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13320_ _18091_/Q _13324_/A _12764_/X vssd1 vssd1 vccd1 vccd1 _13320_/Y sky130_fd_sc_hd__o21ai_1
X_10532_ _10528_/X _10531_/X _10903_/S vssd1 vssd1 vccd1 vccd1 _10532_/X sky130_fd_sc_hd__mux2_1
XFILLER_122_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_210_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_182_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13251_ _13255_/A _18080_/Q vssd1 vssd1 vccd1 vccd1 _13252_/A sky130_fd_sc_hd__and2_1
X_10463_ _09287_/A _09287_/D _09282_/D _09282_/B _10462_/X _10450_/S vssd1 vssd1 vccd1
+ vccd1 _10463_/X sky130_fd_sc_hd__mux4_1
XFILLER_202_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12202_ _11704_/C _12201_/X _12200_/X vssd1 vssd1 vccd1 vccd1 _12202_/Y sky130_fd_sc_hd__o21ai_1
X_13182_ _13186_/A _18049_/Q vssd1 vssd1 vccd1 vccd1 _13183_/A sky130_fd_sc_hd__and2_1
XFILLER_89_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10394_ _10278_/X _10384_/X _10386_/X _10388_/X _10393_/X vssd1 vssd1 vccd1 vccd1
+ _10394_/X sky130_fd_sc_hd__a32o_1
X_12133_ _12133_/A _12133_/B vssd1 vssd1 vccd1 vccd1 _12133_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_150_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17990_ _17990_/CLK _17990_/D vssd1 vssd1 vccd1 vccd1 _17990_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_151_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16941_ _16943_/B _16938_/X _16939_/Y _16940_/X vssd1 vssd1 vccd1 vccd1 _18799_/D
+ sky130_fd_sc_hd__o211a_1
X_12064_ _12066_/A _13420_/A vssd1 vssd1 vccd1 vccd1 _12067_/A sky130_fd_sc_hd__nor2_1
XFILLER_172_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_172_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_1283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11015_ _17999_/Q _17998_/Q vssd1 vssd1 vccd1 vccd1 _11037_/C sky130_fd_sc_hd__nor2_1
XFILLER_42_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16872_ _16874_/B _16869_/X _16870_/Y _16871_/X vssd1 vssd1 vccd1 vccd1 _18784_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_46_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18611_ _18614_/CLK _18611_/D vssd1 vssd1 vccd1 vccd1 _18611_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_49_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15823_ _15823_/A vssd1 vssd1 vccd1 vccd1 _15823_/X sky130_fd_sc_hd__clkbuf_2
XTAP_4040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_219_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18542_ _18542_/CLK _18542_/D vssd1 vssd1 vccd1 vccd1 _18542_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_4084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15754_ _15754_/A _15754_/B vssd1 vssd1 vccd1 vccd1 _15754_/Y sky130_fd_sc_hd__nand2_1
XTAP_4095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINSDIODE2_90 _13752_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12966_ _12966_/A vssd1 vssd1 vccd1 vccd1 _12967_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_166_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14705_ _15145_/A _15145_/B vssd1 vssd1 vccd1 vccd1 _14706_/B sky130_fd_sc_hd__nand2_1
XFILLER_33_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18473_ _18473_/CLK _18473_/D vssd1 vssd1 vccd1 vccd1 _18473_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_3394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11917_ _11917_/A _11917_/B vssd1 vssd1 vccd1 vccd1 _11918_/B sky130_fd_sc_hd__xor2_1
X_15685_ _15982_/A _15696_/B vssd1 vssd1 vccd1 vccd1 _15694_/B sky130_fd_sc_hd__nor2_1
XFILLER_45_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12897_ _12899_/B _12915_/B _12897_/C vssd1 vssd1 vccd1 vccd1 _12898_/A sky130_fd_sc_hd__and3b_1
XTAP_2671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17424_ _18954_/Q _18918_/Q _17427_/S vssd1 vssd1 vccd1 vccd1 _17424_/X sky130_fd_sc_hd__mux2_1
XTAP_2682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14636_ _18251_/Q _14635_/B _14635_/Y _14629_/X vssd1 vssd1 vccd1 vccd1 _18251_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_2693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11848_ _11848_/A _11848_/B vssd1 vssd1 vccd1 vccd1 _11848_/X sky130_fd_sc_hd__or2_1
XFILLER_21_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17355_ _17360_/B _17353_/X _17354_/X _17341_/X vssd1 vssd1 vccd1 vccd1 _18900_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_105_1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14567_ _14690_/B _15172_/A vssd1 vssd1 vccd1 vccd1 _14574_/B sky130_fd_sc_hd__nor2_1
XFILLER_20_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11779_ _11742_/B _11720_/Y _11778_/X vssd1 vssd1 vccd1 vccd1 _11779_/X sky130_fd_sc_hd__o21a_1
XFILLER_53_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16306_ _16305_/B _16304_/X _16305_/Y _16295_/X vssd1 vssd1 vccd1 vccd1 _18647_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_202_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13518_ _13518_/A _13518_/B _13526_/C vssd1 vssd1 vccd1 vccd1 _13552_/B sky130_fd_sc_hd__or3_4
X_17286_ _17464_/A vssd1 vssd1 vccd1 vccd1 _17334_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_201_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14498_ _18223_/Q _14502_/B vssd1 vssd1 vccd1 vccd1 _14499_/A sky130_fd_sc_hd__and2_1
XFILLER_105_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19025_ _19026_/CLK _19025_/D vssd1 vssd1 vccd1 vccd1 _19025_/Q sky130_fd_sc_hd__dfxtp_1
X_16237_ _16248_/A _16678_/B _16272_/C vssd1 vssd1 vccd1 vccd1 _16237_/X sky130_fd_sc_hd__or3_1
XFILLER_173_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13449_ _11720_/B _13448_/Y _11333_/Y _11586_/A vssd1 vssd1 vccd1 vccd1 _13449_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_220_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_75_wb_clk_i clkbuf_5_21_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18682_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_103_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16168_ _16181_/A _16759_/B _16181_/C vssd1 vssd1 vccd1 vccd1 _16168_/X sky130_fd_sc_hd__or3_1
XFILLER_154_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_216_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15119_ _15118_/B _15117_/X _15118_/Y _15103_/X vssd1 vssd1 vccd1 vccd1 _18368_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_142_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16099_ _16850_/A vssd1 vssd1 vccd1 vccd1 _16701_/A sky130_fd_sc_hd__buf_8
X_08990_ _08991_/A vssd1 vssd1 vccd1 vccd1 _08990_/Y sky130_fd_sc_hd__inv_2
XFILLER_69_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_214_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_205_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_96_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_217_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_214_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09611_ _09611_/A _09611_/B vssd1 vssd1 vccd1 vccd1 _10110_/A sky130_fd_sc_hd__xnor2_4
XFILLER_112_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18809_ _18809_/CLK _18809_/D vssd1 vssd1 vccd1 vccd1 _18809_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_28_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_216_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09542_ _10007_/B vssd1 vssd1 vccd1 vccd1 _12066_/A sky130_fd_sc_hd__buf_2
XFILLER_209_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09473_ _09474_/A _09457_/B _18142_/D vssd1 vssd1 vccd1 vccd1 _18139_/D sky130_fd_sc_hd__a21o_1
XFILLER_24_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_225_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_221_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_212_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_212_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_192_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_164_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_182_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19086__57 vssd1 vssd1 vccd1 vccd1 _19086__57/HI _19194_/A sky130_fd_sc_hd__conb_1
XFILLER_191_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09809_ _09810_/B _09810_/C _09810_/A vssd1 vssd1 vccd1 vccd1 _12106_/A sky130_fd_sc_hd__a21oi_1
XFILLER_207_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_219_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_216_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12820_ _17933_/Q _12795_/Y _12798_/Y _17937_/Q vssd1 vssd1 vccd1 vccd1 _12820_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_75_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12751_ _18025_/Q _18024_/Q _18027_/Q _18026_/Q vssd1 vssd1 vccd1 vccd1 _12752_/C
+ sky130_fd_sc_hd__and4_1
XTAP_1211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_216_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11702_ _11704_/A _11390_/X _11700_/Y _11848_/A vssd1 vssd1 vccd1 vccd1 _11702_/X
+ sky130_fd_sc_hd__a31o_1
XTAP_1244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15470_ _18447_/Q _15473_/B _15469_/X _15452_/X vssd1 vssd1 vccd1 vccd1 _18447_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_1255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12682_ _17937_/Q vssd1 vssd1 vccd1 vccd1 _12707_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_128_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14421_ _14421_/A vssd1 vssd1 vccd1 vccd1 _14452_/A sky130_fd_sc_hd__buf_2
XFILLER_70_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11633_ _11770_/C _11633_/B vssd1 vssd1 vccd1 vccd1 _11757_/A sky130_fd_sc_hd__and2_1
XFILLER_230_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17140_ _17197_/A vssd1 vssd1 vccd1 vccd1 _17140_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_211_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14352_ _18182_/Q vssd1 vssd1 vccd1 vccd1 _17575_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_196_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11564_ _11549_/X _11565_/B _11560_/X _11563_/X vssd1 vssd1 vccd1 vccd1 _11564_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_168_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13303_ _13303_/A _13303_/B _13303_/C vssd1 vssd1 vccd1 vccd1 _13304_/B sky130_fd_sc_hd__or3_1
X_17071_ _18867_/Q _18831_/Q _17074_/S vssd1 vssd1 vccd1 vccd1 _17071_/X sky130_fd_sc_hd__mux2_1
X_10515_ _14307_/A _10939_/C _10515_/C vssd1 vssd1 vccd1 vccd1 _10515_/X sky130_fd_sc_hd__and3_1
XFILLER_144_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11495_ _11261_/X _11495_/B _13444_/A _11495_/D vssd1 vssd1 vccd1 vccd1 _11501_/B
+ sky130_fd_sc_hd__and4b_1
XFILLER_6_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14283_ _14283_/A vssd1 vssd1 vccd1 vccd1 _14283_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_183_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16022_ _16027_/B _16020_/X _16021_/X _16008_/X vssd1 vssd1 vccd1 vccd1 _18582_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_171_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13234_ _13234_/A vssd1 vssd1 vccd1 vccd1 _18071_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_87_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10446_ _09253_/A _09243_/D _10503_/S vssd1 vssd1 vccd1 vccd1 _10446_/X sky130_fd_sc_hd__mux2_1
XFILLER_171_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_226_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_174_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10377_ _09327_/A _10316_/S _10376_/X _09948_/A vssd1 vssd1 vccd1 vccd1 _10377_/X
+ sky130_fd_sc_hd__o211a_1
X_13165_ _13165_/A vssd1 vssd1 vccd1 vccd1 _18040_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_100_1288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_1367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12116_ _17977_/Q _12116_/B vssd1 vssd1 vccd1 vccd1 _12117_/B sky130_fd_sc_hd__xnor2_1
X_13096_ _13096_/A vssd1 vssd1 vccd1 vccd1 _18009_/D sky130_fd_sc_hd__clkbuf_1
X_17973_ _17990_/CLK _17973_/D vssd1 vssd1 vccd1 vccd1 _17973_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_111_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_215_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16924_ _16930_/B _16921_/X _16923_/X _16917_/X vssd1 vssd1 vccd1 vccd1 _18795_/D
+ sky130_fd_sc_hd__o211a_1
X_12047_ _12047_/A _12133_/B vssd1 vssd1 vccd1 vccd1 _12054_/B sky130_fd_sc_hd__nor2_1
XFILLER_78_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_193_wb_clk_i clkbuf_5_9_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18209_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_16855_ _16860_/B _16852_/X _16854_/X _16848_/X vssd1 vssd1 vccd1 vccd1 _18780_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_225_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15806_ _15818_/A _15806_/B vssd1 vssd1 vccd1 vccd1 _15806_/Y sky130_fd_sc_hd__nand2_1
Xclkbuf_leaf_122_wb_clk_i clkbuf_5_25_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18432_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_81_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16786_ _16792_/B _16784_/X _16785_/X _16781_/X vssd1 vssd1 vccd1 vccd1 _18765_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_225_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13998_ _18562_/Q _13749_/A _13994_/X _13997_/X vssd1 vssd1 vccd1 vccd1 _13998_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18525_ _18572_/CLK _18525_/D vssd1 vssd1 vccd1 vccd1 _18525_/Q sky130_fd_sc_hd__dfxtp_4
X_15737_ _18550_/Q _18514_/Q _15753_/S vssd1 vssd1 vccd1 vccd1 _15737_/X sky130_fd_sc_hd__mux2_1
XTAP_3180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12949_ _12760_/A _12947_/X _12948_/X _12928_/X vssd1 vssd1 vccd1 vccd1 _12949_/Y
+ sky130_fd_sc_hd__o31ai_4
XFILLER_222_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18456_ _18458_/CLK _18456_/D vssd1 vssd1 vccd1 vccd1 _18456_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_222_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15668_ _15717_/A vssd1 vssd1 vccd1 vccd1 _15693_/S sky130_fd_sc_hd__clkbuf_2
XTAP_2490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_178_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17407_ _17468_/A vssd1 vssd1 vccd1 vccd1 _17456_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_222_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14619_ _14360_/X _14608_/X _14612_/X _14617_/Y _14618_/X vssd1 vssd1 vccd1 vccd1
+ _18248_/D sky130_fd_sc_hd__o311a_1
XFILLER_60_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18387_ _18387_/CLK _18387_/D vssd1 vssd1 vccd1 vccd1 _18387_/Q sky130_fd_sc_hd__dfxtp_2
X_15599_ _15613_/A _16043_/B _15599_/C vssd1 vssd1 vccd1 vccd1 _15599_/X sky130_fd_sc_hd__or3_1
XFILLER_159_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_193_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_159_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17338_ _17480_/A _17351_/B vssd1 vssd1 vccd1 vccd1 _17349_/B sky130_fd_sc_hd__nor2_1
XFILLER_140_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17269_ _17331_/A vssd1 vssd1 vccd1 vccd1 _17397_/B sky130_fd_sc_hd__buf_2
XFILLER_179_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19008_ _19009_/CLK _19008_/D vssd1 vssd1 vccd1 vccd1 _19008_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_106_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_216_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08973_ input1/X vssd1 vssd1 vccd1 vccd1 _08998_/A sky130_fd_sc_hd__buf_4
XFILLER_103_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_216_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_151_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_1295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09525_ _14199_/A vssd1 vssd1 vccd1 vccd1 _14299_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_227_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_213_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_225_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_3_5_0_wb_clk_i clkbuf_3_5_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_5_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_2
XPHY_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_227_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09456_ _09463_/A _09475_/B vssd1 vssd1 vccd1 vccd1 _09457_/B sky130_fd_sc_hd__or2_2
XFILLER_212_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_212_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_197_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09387_ _09387_/A _09387_/B _09387_/C vssd1 vssd1 vccd1 vccd1 _09450_/A sky130_fd_sc_hd__and3_2
XFILLER_177_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_1277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10300_ _09214_/A _09219_/C _09219_/D _09209_/B _10376_/B _09953_/A vssd1 vssd1 vccd1
+ vccd1 _10300_/X sky130_fd_sc_hd__mux4_1
XFILLER_158_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11280_ _11590_/B _11334_/B vssd1 vssd1 vccd1 vccd1 _11280_/Y sky130_fd_sc_hd__nor2_1
XFILLER_146_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10231_ _10489_/S vssd1 vssd1 vccd1 vccd1 _10231_/X sky130_fd_sc_hd__buf_4
XFILLER_106_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10162_ _10162_/A _10168_/B vssd1 vssd1 vccd1 vccd1 _10178_/B sky130_fd_sc_hd__xnor2_2
XFILLER_133_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14970_ _18368_/Q _18332_/Q _14974_/S vssd1 vssd1 vccd1 vccd1 _14970_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10093_ _09657_/A _10940_/A _10082_/X _10092_/Y vssd1 vssd1 vccd1 vccd1 _10093_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_43_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13921_ _18751_/Q _13568_/A _13919_/X _13920_/X vssd1 vssd1 vccd1 vccd1 _13921_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_48_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16640_ _16648_/B _16637_/X _16638_/X _16639_/X vssd1 vssd1 vccd1 vccd1 _18729_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_130_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13852_ _18718_/Q _13523_/A _13598_/X _18700_/Q vssd1 vssd1 vccd1 vccd1 _13852_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_47_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_216_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12803_ _17947_/Q vssd1 vssd1 vccd1 vccd1 _12846_/A sky130_fd_sc_hd__inv_2
X_16571_ _18748_/Q _18712_/Q _16598_/S vssd1 vssd1 vccd1 vccd1 _16571_/X sky130_fd_sc_hd__mux2_1
X_13783_ _18426_/Q _13580_/A _13734_/X _18420_/Q _13782_/X vssd1 vssd1 vccd1 vccd1
+ _13783_/X sky130_fd_sc_hd__a221o_1
XFILLER_128_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10995_ _18995_/Q _09523_/X _10977_/A _10982_/A _14267_/A vssd1 vssd1 vccd1 vccd1
+ _18995_/D sky130_fd_sc_hd__a32o_1
X_18310_ _18324_/CLK _18310_/D vssd1 vssd1 vccd1 vccd1 _18310_/Q sky130_fd_sc_hd__dfxtp_4
X_15522_ _15525_/B _15519_/X _15521_/Y _15516_/X vssd1 vssd1 vccd1 vccd1 _18460_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_167_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12734_ _19020_/Q _19019_/Q _19022_/Q _19021_/Q vssd1 vssd1 vccd1 vccd1 _12736_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_215_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_231_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18241_ _18245_/CLK _18241_/D vssd1 vssd1 vccd1 vccd1 _18241_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_128_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15453_ _15460_/B _15449_/X _15451_/X _15452_/X vssd1 vssd1 vccd1 vccd1 _18444_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_1085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12665_ _12665_/A _12665_/B vssd1 vssd1 vccd1 vccd1 _12665_/Y sky130_fd_sc_hd__nand2_1
XFILLER_231_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14404_ _14404_/A vssd1 vssd1 vccd1 vccd1 _14404_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_198_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11616_ _11615_/A _12233_/A _11623_/B _11614_/Y _11615_/Y vssd1 vssd1 vccd1 vccd1
+ _11616_/Y sky130_fd_sc_hd__o311ai_1
XFILLER_15_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18172_ _18184_/CLK _18172_/D vssd1 vssd1 vccd1 vccd1 _18172_/Q sky130_fd_sc_hd__dfxtp_2
X_15384_ _18466_/Q _18430_/Q _15388_/S vssd1 vssd1 vccd1 vccd1 _15384_/X sky130_fd_sc_hd__mux2_1
X_12596_ _17927_/Q _12597_/B vssd1 vssd1 vccd1 vccd1 _12598_/A sky130_fd_sc_hd__and2_1
XFILLER_129_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17123_ _17184_/A vssd1 vssd1 vccd1 vccd1 _17254_/B sky130_fd_sc_hd__buf_2
XFILLER_15_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14335_ _14470_/A _14335_/B vssd1 vssd1 vccd1 vccd1 _14335_/X sky130_fd_sc_hd__or2_1
XFILLER_102_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11547_ _11621_/B _11547_/B vssd1 vssd1 vccd1 vccd1 _11547_/Y sky130_fd_sc_hd__nor2_1
XFILLER_184_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17054_ _17056_/B _17052_/X _17053_/Y _17040_/X vssd1 vssd1 vccd1 vccd1 _18826_/D
+ sky130_fd_sc_hd__o211a_1
X_14266_ _11920_/B _14205_/X _14265_/X vssd1 vssd1 vccd1 vccd1 _14266_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_171_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11478_ _11478_/A _11478_/B vssd1 vssd1 vccd1 vccd1 _11478_/Y sky130_fd_sc_hd__nand2_1
XFILLER_109_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16005_ _16005_/A _16041_/B vssd1 vssd1 vccd1 vccd1 _16017_/B sky130_fd_sc_hd__nor2_2
X_13217_ _13217_/A vssd1 vssd1 vccd1 vccd1 _18063_/D sky130_fd_sc_hd__clkbuf_1
X_10429_ _10494_/A vssd1 vssd1 vccd1 vccd1 _10429_/X sky130_fd_sc_hd__clkbuf_8
XFILLER_171_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14197_ _18218_/Q _18217_/Q _18216_/Q _18215_/Q vssd1 vssd1 vccd1 vccd1 _14216_/A
+ sky130_fd_sc_hd__or4_2
XFILLER_100_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_1262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_125_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13148_ _13148_/A vssd1 vssd1 vccd1 vccd1 _18032_/D sky130_fd_sc_hd__clkbuf_1
XTAP_825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13079_ _13076_/X _13077_/X _13078_/Y vssd1 vssd1 vccd1 vccd1 _18002_/D sky130_fd_sc_hd__o21a_1
X_17956_ _17959_/CLK _17956_/D vssd1 vssd1 vccd1 vccd1 _17956_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16907_ _16928_/A vssd1 vssd1 vccd1 vccd1 _16925_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_22_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17887_ _17890_/CLK _17887_/D vssd1 vssd1 vccd1 vccd1 _17887_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_65_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16838_ _18813_/Q _18777_/Q _16842_/S vssd1 vssd1 vccd1 vccd1 _16838_/X sky130_fd_sc_hd__mux2_1
XFILLER_4_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16769_ _16815_/A _16769_/B vssd1 vssd1 vccd1 vccd1 _16769_/Y sky130_fd_sc_hd__nand2_1
XFILLER_65_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_202_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09310_ _18467_/Q _18466_/Q _18465_/Q vssd1 vssd1 vccd1 vccd1 _09314_/A sky130_fd_sc_hd__or3_4
X_18508_ _18511_/CLK _18508_/D vssd1 vssd1 vccd1 vccd1 _18508_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_55_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_222_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09241_ _18899_/Q _18898_/Q _18897_/Q vssd1 vssd1 vccd1 vccd1 _09243_/C sky130_fd_sc_hd__or3_4
X_18439_ _18443_/CLK _18439_/D vssd1 vssd1 vccd1 vccd1 _18439_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_146_1277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_222_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_90_wb_clk_i clkbuf_5_20_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18662_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_194_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09172_ _18611_/Q _18610_/Q _18609_/Q vssd1 vssd1 vccd1 vccd1 _09176_/A sky130_fd_sc_hd__or3_4
XFILLER_193_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_115_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_6008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_6019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_1264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19056__27 vssd1 vssd1 vccd1 vccd1 _19056__27/HI _19150_/A sky130_fd_sc_hd__conb_1
XFILLER_103_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08956_ _08960_/A vssd1 vssd1 vccd1 vccd1 _08956_/Y sky130_fd_sc_hd__inv_2
XFILLER_131_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_229_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_116_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_229_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_217_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_229_1319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09508_ _14297_/A _17704_/A vssd1 vssd1 vccd1 vccd1 _09518_/B sky130_fd_sc_hd__or2_1
XPHY_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10780_ _09332_/B _09327_/B _09337_/C _09327_/C _10687_/A _10743_/A vssd1 vssd1 vccd1
+ vccd1 _10780_/X sky130_fd_sc_hd__mux4_2
XFILLER_213_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_1366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09439_ _09439_/A vssd1 vssd1 vccd1 vccd1 _18134_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_38_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_212_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12450_ _17903_/Q _12450_/B vssd1 vssd1 vccd1 vccd1 _12451_/B sky130_fd_sc_hd__or2_1
XFILLER_40_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_227_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11401_ _11442_/A _11442_/B vssd1 vssd1 vccd1 vccd1 _11652_/A sky130_fd_sc_hd__and2_1
XFILLER_165_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12381_ _18105_/Q _12381_/B vssd1 vssd1 vccd1 vccd1 _12384_/B sky130_fd_sc_hd__and2b_1
XFILLER_193_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14120_ _18947_/Q _13838_/X _14015_/X _18950_/Q _14119_/X vssd1 vssd1 vccd1 vccd1
+ _14120_/X sky130_fd_sc_hd__a221o_1
X_11332_ _11330_/Y _17875_/Q _11331_/X _17877_/Q vssd1 vssd1 vccd1 vccd1 _11332_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_21_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14051_ _18506_/Q _13561_/A _13492_/A _18497_/Q vssd1 vssd1 vccd1 vccd1 _14051_/X
+ sky130_fd_sc_hd__a22o_1
X_11263_ _17803_/Q _12036_/B vssd1 vssd1 vccd1 vccd1 _12037_/A sky130_fd_sc_hd__or2_2
XFILLER_4_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13002_ _17990_/Q _12955_/X _13001_/Y _12721_/X _13007_/B vssd1 vssd1 vccd1 vccd1
+ _13002_/X sky130_fd_sc_hd__a221o_1
XFILLER_106_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_122_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10214_ _10218_/A _10218_/B vssd1 vssd1 vccd1 vccd1 _10215_/B sky130_fd_sc_hd__xnor2_2
XFILLER_121_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11194_ _11210_/A _11194_/B vssd1 vssd1 vccd1 vccd1 _11195_/A sky130_fd_sc_hd__and2_1
XFILLER_161_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17810_ _18989_/CLK _17810_/D vssd1 vssd1 vccd1 vccd1 _17810_/Q sky130_fd_sc_hd__dfxtp_1
X_10145_ _10146_/A _10146_/B vssd1 vssd1 vccd1 vccd1 _10147_/A sky130_fd_sc_hd__nor2_1
X_18790_ _18826_/CLK _18790_/D vssd1 vssd1 vccd1 vccd1 _18790_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_5830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17741_ _17745_/A _19015_/Q vssd1 vssd1 vccd1 vccd1 _17742_/A sky130_fd_sc_hd__and2_1
XFILLER_94_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14953_ _14975_/A _15243_/B _14965_/C vssd1 vssd1 vccd1 vccd1 _14953_/X sky130_fd_sc_hd__or3_1
X_10076_ _10074_/X _10075_/X _10076_/S vssd1 vssd1 vccd1 vccd1 _10076_/X sky130_fd_sc_hd__mux2_1
XFILLER_43_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13904_ _18544_/Q _13731_/A _13630_/A _18520_/Q _13903_/X vssd1 vssd1 vccd1 vccd1
+ _13904_/X sky130_fd_sc_hd__a221o_1
X_17672_ _17681_/A _17672_/B vssd1 vssd1 vccd1 vccd1 _17673_/A sky130_fd_sc_hd__and2_1
XFILLER_78_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14884_ _14944_/A vssd1 vssd1 vccd1 vccd1 _14932_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_63_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16623_ _16634_/A _16623_/B vssd1 vssd1 vccd1 vccd1 _16623_/Y sky130_fd_sc_hd__nand2_1
X_19070__41 vssd1 vssd1 vccd1 vccd1 _19070__41/HI _19164_/A sky130_fd_sc_hd__conb_1
X_13835_ _18676_/Q _13493_/X _13500_/X _18691_/Q vssd1 vssd1 vccd1 vccd1 _13835_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_90_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_204 _12346_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINSDIODE2_215 _13715_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_226 _15175_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16554_ _18744_/Q _18708_/Q _16565_/S vssd1 vssd1 vccd1 vccd1 _16554_/X sky130_fd_sc_hd__mux2_1
XPHY_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XINSDIODE2_237 _17814_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13766_ _13766_/A vssd1 vssd1 vccd1 vccd1 _13766_/X sky130_fd_sc_hd__buf_4
XINSDIODE2_248 _09098_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_188_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_259 _13834_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10978_ _14299_/A vssd1 vssd1 vccd1 vccd1 _14272_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_206_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_1327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15505_ _15551_/A _15946_/B _15515_/C vssd1 vssd1 vccd1 vccd1 _15505_/X sky130_fd_sc_hd__or3_1
XFILLER_231_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12717_ _12951_/A vssd1 vssd1 vccd1 vccd1 _12962_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_203_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16485_ _16487_/B _16483_/X _16484_/Y _16477_/X vssd1 vssd1 vccd1 vccd1 _18691_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_43_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13697_ _13697_/A vssd1 vssd1 vccd1 vccd1 _13698_/A sky130_fd_sc_hd__buf_2
XFILLER_30_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_206_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18224_ _18224_/CLK _18224_/D vssd1 vssd1 vccd1 vccd1 _18224_/Q sky130_fd_sc_hd__dfxtp_1
X_15436_ _15562_/A vssd1 vssd1 vccd1 vccd1 _15492_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_188_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12648_ _12640_/A _12640_/B _12638_/A vssd1 vssd1 vccd1 vccd1 _12649_/B sky130_fd_sc_hd__a21o_1
XFILLER_15_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18155_ _18157_/CLK _18155_/D vssd1 vssd1 vccd1 vccd1 _18155_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15367_ _15366_/B _15365_/X _15366_/Y _15363_/X vssd1 vssd1 vccd1 vccd1 _18425_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_200_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12579_ _17925_/Q _17922_/Q vssd1 vssd1 vccd1 vccd1 _12580_/A sky130_fd_sc_hd__xnor2_1
XFILLER_156_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17106_ _17105_/B _17103_/X _17105_/Y _17096_/X vssd1 vssd1 vccd1 vccd1 _18839_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_89_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14318_ _12101_/A _14188_/A _14307_/B _10939_/C _14317_/Y vssd1 vssd1 vccd1 vccd1
+ _14318_/X sky130_fd_sc_hd__o221a_1
XFILLER_102_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18086_ _18087_/CLK _18086_/D vssd1 vssd1 vccd1 vccd1 _18086_/Q sky130_fd_sc_hd__dfxtp_1
X_15298_ _15448_/B vssd1 vssd1 vccd1 vccd1 _15358_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_183_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17037_ _17037_/A _17109_/C vssd1 vssd1 vccd1 vccd1 _17046_/B sky130_fd_sc_hd__nor2_2
XFILLER_176_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14249_ _14248_/X _09981_/X _14260_/A vssd1 vssd1 vccd1 vccd1 _14249_/X sky130_fd_sc_hd__mux2_1
XFILLER_217_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_139_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09790_ _09891_/A _09891_/B vssd1 vssd1 vccd1 vccd1 _09790_/X sky130_fd_sc_hd__and2b_1
XTAP_666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18988_ _18988_/CLK _18988_/D vssd1 vssd1 vccd1 vccd1 _18988_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17939_ _17939_/CLK _17939_/D vssd1 vssd1 vccd1 vccd1 _17939_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_66_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_226_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_213_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_227_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_227_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_1238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_226_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_224_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_210_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09224_ _18923_/Q _18922_/Q _18921_/Q vssd1 vssd1 vccd1 vccd1 _09227_/B sky130_fd_sc_hd__or3_4
XFILLER_33_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_1361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09155_ _09431_/A _09429_/A vssd1 vssd1 vccd1 vccd1 _09222_/A sky130_fd_sc_hd__nor2_1
XFILLER_175_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09086_ _09086_/A vssd1 vssd1 vccd1 vccd1 _19181_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_120_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_225_wb_clk_i _17864_/CLK vssd1 vssd1 vccd1 vccd1 _17895_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_190_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_5_26_0_wb_clk_i clkbuf_5_27_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_5_26_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_118_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09988_ _09153_/A _09143_/B _09148_/C _10722_/A _10955_/S _09987_/X vssd1 vssd1 vccd1
+ vccd1 _09988_/X sky130_fd_sc_hd__mux4_1
XFILLER_130_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08939_ _08941_/A vssd1 vssd1 vccd1 vccd1 _08939_/Y sky130_fd_sc_hd__inv_2
XTAP_4425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_218_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11950_ _11939_/X _11944_/X _12049_/A vssd1 vssd1 vccd1 vccd1 _12028_/D sky130_fd_sc_hd__a21oi_4
XFILLER_229_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10901_ _09413_/C _09418_/B _09408_/A _09408_/B _10542_/X _10518_/X vssd1 vssd1 vccd1
+ vccd1 _10901_/X sky130_fd_sc_hd__mux4_2
XTAP_3768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11881_ _13210_/A vssd1 vssd1 vccd1 vccd1 _12207_/A sky130_fd_sc_hd__buf_4
XFILLER_72_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13620_ _18477_/Q _13617_/X _13619_/X _18453_/Q vssd1 vssd1 vccd1 vccd1 _13620_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_199_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10832_ _10700_/S _10838_/B _10823_/X _10828_/X _10831_/X vssd1 vssd1 vccd1 vccd1
+ _10833_/C sky130_fd_sc_hd__o311a_1
XFILLER_25_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_213_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13551_ _13837_/A vssd1 vssd1 vccd1 vccd1 _13551_/X sky130_fd_sc_hd__buf_2
XFILLER_38_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_198_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10763_ _09186_/B _09181_/C _10763_/S vssd1 vssd1 vccd1 vccd1 _10764_/B sky130_fd_sc_hd__mux2_1
XFILLER_41_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12502_ _17911_/Q _12501_/X _12472_/A vssd1 vssd1 vccd1 vccd1 _12502_/Y sky130_fd_sc_hd__o21ai_1
X_16270_ _16714_/A _16307_/B vssd1 vssd1 vccd1 vccd1 _16285_/B sky130_fd_sc_hd__nor2_1
X_13482_ _17848_/Q _13464_/X _13465_/A vssd1 vssd1 vccd1 vccd1 _13483_/B sky130_fd_sc_hd__a21oi_1
X_10694_ _09198_/A _09193_/A _09203_/B _10293_/A _10693_/X _10680_/A vssd1 vssd1 vccd1
+ vccd1 _10694_/X sky130_fd_sc_hd__mux4_1
XFILLER_125_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15221_ _15227_/B _15219_/X _15220_/X _15208_/X vssd1 vssd1 vccd1 vccd1 _18393_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_185_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12433_ _12433_/A vssd1 vssd1 vccd1 vccd1 _17900_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_12_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15152_ _15178_/A _15154_/B vssd1 vssd1 vccd1 vccd1 _15152_/Y sky130_fd_sc_hd__nand2_1
XFILLER_154_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12364_ _18989_/Q vssd1 vssd1 vccd1 vccd1 _12373_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_148_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14103_ _18662_/Q _14015_/A _14027_/A _18653_/Q _14102_/X vssd1 vssd1 vccd1 vccd1
+ _14103_/X sky130_fd_sc_hd__a221o_2
XFILLER_181_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11315_ _11368_/B _11315_/B _13443_/A _11368_/A vssd1 vssd1 vccd1 vccd1 _11316_/B
+ sky130_fd_sc_hd__and4b_1
X_15083_ _15083_/A vssd1 vssd1 vccd1 vccd1 _15083_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_153_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12295_ _17873_/Q _12287_/Y _12313_/B vssd1 vssd1 vccd1 vccd1 _17873_/D sky130_fd_sc_hd__o21a_1
X_14034_ _18239_/Q _13619_/X _14029_/X _14033_/X vssd1 vssd1 vccd1 vccd1 _14034_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_49_1262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18911_ _18927_/CLK _18911_/D vssd1 vssd1 vccd1 vccd1 _18911_/Q sky130_fd_sc_hd__dfxtp_2
X_11246_ _11245_/A _11245_/B _11245_/Y _11221_/X vssd1 vssd1 vccd1 vccd1 _17824_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_180_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18842_ _18845_/CLK _18842_/D vssd1 vssd1 vccd1 vccd1 _18842_/Q sky130_fd_sc_hd__dfxtp_1
X_11177_ _17806_/Q _11177_/B vssd1 vssd1 vccd1 vccd1 _11178_/C sky130_fd_sc_hd__or2_1
XFILLER_110_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_212_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10128_ _18127_/Q vssd1 vssd1 vccd1 vccd1 _10159_/A sky130_fd_sc_hd__clkbuf_4
X_15985_ _15991_/B _15983_/X _15984_/X _15972_/X vssd1 vssd1 vccd1 vccd1 _18573_/D
+ sky130_fd_sc_hd__o211a_1
X_18773_ _18773_/CLK _18773_/D vssd1 vssd1 vccd1 vccd1 _18773_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_5660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14936_ _14935_/B _14934_/X _14935_/Y _14922_/X vssd1 vssd1 vccd1 vccd1 _18323_/D
+ sky130_fd_sc_hd__o211a_1
X_10059_ _09209_/A _09219_/B _09214_/D _09214_/B _09703_/A _09709_/A vssd1 vssd1 vccd1
+ vccd1 _10059_/X sky130_fd_sc_hd__mux4_1
X_17724_ _17724_/A vssd1 vssd1 vccd1 vccd1 _19006_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_76_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_212_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_208_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_29_wb_clk_i clkbuf_5_5_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18914_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_4992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14867_ _18342_/Q _18306_/Q _14883_/S vssd1 vssd1 vccd1 vccd1 _14867_/X sky130_fd_sc_hd__mux2_1
X_17655_ _17641_/X _17649_/Y _17654_/X _17650_/Y _18976_/Q vssd1 vssd1 vccd1 vccd1
+ _17656_/B sky130_fd_sc_hd__a32o_1
XFILLER_21_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16606_ _16611_/B _16604_/X _16605_/X _16600_/X vssd1 vssd1 vccd1 vccd1 _18720_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_51_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13818_ _18921_/Q _13733_/A _13814_/X _13817_/X vssd1 vssd1 vccd1 vccd1 _13818_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_1_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17586_ _17571_/X _17576_/Y _17582_/X _17577_/Y _18959_/Q vssd1 vssd1 vccd1 vccd1
+ _17587_/B sky130_fd_sc_hd__a32o_1
XFILLER_91_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14798_ _15207_/A vssd1 vssd1 vccd1 vccd1 _14881_/A sky130_fd_sc_hd__buf_2
XFILLER_189_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16537_ _18740_/Q _18704_/Q _16546_/S vssd1 vssd1 vccd1 vccd1 _16537_/X sky130_fd_sc_hd__mux2_1
X_13749_ _13749_/A vssd1 vssd1 vccd1 vccd1 _13749_/X sky130_fd_sc_hd__buf_6
XFILLER_92_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16468_ _16491_/A _16759_/B _16481_/C vssd1 vssd1 vccd1 vccd1 _16468_/X sky130_fd_sc_hd__or3_1
XFILLER_143_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15419_ _16935_/A vssd1 vssd1 vccd1 vccd1 _16019_/A sky130_fd_sc_hd__clkbuf_4
X_18207_ _18992_/CLK _18207_/D vssd1 vssd1 vccd1 vccd1 _18207_/Q sky130_fd_sc_hd__dfxtp_1
X_19187_ _19187_/A _09003_/Y vssd1 vssd1 vccd1 vccd1 io_out[25] sky130_fd_sc_hd__ebufn_8
X_16399_ _16407_/B _16396_/X _16397_/X _16398_/X vssd1 vssd1 vccd1 vccd1 _18669_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_191_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18138_ _18140_/CLK _18138_/D vssd1 vssd1 vccd1 vccd1 _18138_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_163_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18069_ _18069_/CLK _18069_/D vssd1 vssd1 vccd1 vccd1 _18069_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_208_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09911_ _09962_/A vssd1 vssd1 vccd1 vccd1 _09953_/A sky130_fd_sc_hd__buf_4
XFILLER_208_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09842_ _12109_/B _09842_/B vssd1 vssd1 vccd1 vccd1 _09843_/B sky130_fd_sc_hd__xnor2_1
XFILLER_112_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_224_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09773_ _18101_/Q vssd1 vssd1 vccd1 vccd1 _09918_/A sky130_fd_sc_hd__inv_2
XTAP_496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_230_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_224_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_227_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_230_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_226_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_215_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_214_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_224_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_223_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_224_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09207_ _18677_/Q _18676_/Q _18675_/Q vssd1 vssd1 vccd1 vccd1 _09209_/C sky130_fd_sc_hd__or3_4
XFILLER_194_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09138_ _09138_/A _09138_/B vssd1 vssd1 vccd1 vccd1 _09431_/A sky130_fd_sc_hd__or2_1
XFILLER_68_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_123_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09069_ _09072_/A _09069_/B _17828_/Q vssd1 vssd1 vccd1 vccd1 _09070_/A sky130_fd_sc_hd__and3_1
XFILLER_118_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11100_ _17795_/Q vssd1 vssd1 vccd1 vccd1 _11586_/A sky130_fd_sc_hd__buf_2
XFILLER_118_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12080_ _12079_/Y _09684_/A _12080_/S vssd1 vssd1 vccd1 vccd1 _12080_/X sky130_fd_sc_hd__mux2_1
XFILLER_1_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_104_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11031_ _11031_/A _13337_/A vssd1 vssd1 vccd1 vccd1 _11031_/X sky130_fd_sc_hd__or2_2
XFILLER_134_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15770_ _18521_/Q _15769_/B _15769_/Y _15763_/X vssd1 vssd1 vccd1 vccd1 _18521_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_4255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12982_ _12982_/A _12982_/B vssd1 vssd1 vccd1 vccd1 _12983_/B sky130_fd_sc_hd__xnor2_1
XFILLER_57_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14721_ _14812_/A vssd1 vssd1 vccd1 vccd1 _14736_/S sky130_fd_sc_hd__clkbuf_2
XTAP_3543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_218_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11933_ _11964_/A _11979_/A _11983_/B _11983_/A vssd1 vssd1 vccd1 vccd1 _12007_/B
+ sky130_fd_sc_hd__o211a_2
XFILLER_79_1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19040__11 vssd1 vssd1 vccd1 vccd1 _19040__11/HI _19134_/A sky130_fd_sc_hd__conb_1
XFILLER_75_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17440_ _17453_/A _17444_/B vssd1 vssd1 vccd1 vccd1 _17440_/Y sky130_fd_sc_hd__nand2_1
XTAP_2842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14652_ _16919_/A vssd1 vssd1 vccd1 vccd1 _16922_/A sky130_fd_sc_hd__buf_4
XTAP_3598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11864_ _18157_/Q _11813_/Y _11861_/X _11863_/X vssd1 vssd1 vccd1 vccd1 _17828_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_73_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13603_ _18825_/Q _13525_/A _13546_/X _18813_/Q vssd1 vssd1 vccd1 vccd1 _13603_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_2886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17371_ _18941_/Q _18905_/Q _17386_/S vssd1 vssd1 vccd1 vccd1 _17371_/X sky130_fd_sc_hd__mux2_1
XTAP_2897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10815_ _10702_/A _10812_/X _10814_/X _10805_/A vssd1 vssd1 vccd1 vccd1 _10815_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_214_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14583_ _16853_/A vssd1 vssd1 vccd1 vccd1 _15186_/B sky130_fd_sc_hd__buf_8
X_11795_ _11795_/A _11795_/B vssd1 vssd1 vccd1 vccd1 _11797_/B sky130_fd_sc_hd__xnor2_1
XFILLER_129_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16322_ _16371_/A _16759_/B _16333_/C vssd1 vssd1 vccd1 vccd1 _16322_/X sky130_fd_sc_hd__or3_1
XFILLER_14_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13534_ _13724_/A vssd1 vssd1 vccd1 vccd1 _13535_/A sky130_fd_sc_hd__buf_2
XFILLER_201_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10746_ _09119_/A _09109_/D _10810_/S vssd1 vssd1 vccd1 vccd1 _10747_/B sky130_fd_sc_hd__mux2_1
XFILLER_14_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16253_ _16256_/B _16250_/X _16251_/Y _16252_/X vssd1 vssd1 vccd1 vccd1 _18634_/D
+ sky130_fd_sc_hd__o211a_1
Xclkbuf_leaf_147_wb_clk_i clkbuf_5_26_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18299_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_16_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13465_ _13465_/A vssd1 vssd1 vccd1 vccd1 _13465_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_51_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10677_ _10833_/A vssd1 vssd1 vccd1 vccd1 _10910_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_103_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15204_ _15206_/B _15202_/X _15203_/Y _15187_/X vssd1 vssd1 vccd1 vccd1 _18388_/D
+ sky130_fd_sc_hd__o211a_1
X_12416_ _12416_/A vssd1 vssd1 vccd1 vccd1 _17898_/D sky130_fd_sc_hd__clkbuf_1
X_16184_ _16199_/A _16188_/B vssd1 vssd1 vccd1 vccd1 _16184_/Y sky130_fd_sc_hd__nand2_1
XFILLER_173_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13396_ _18123_/Q _11021_/X _13342_/X _13395_/X vssd1 vssd1 vccd1 vccd1 _18123_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_182_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_177_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15135_ _18408_/Q _18372_/Q _15141_/S vssd1 vssd1 vccd1 vccd1 _15135_/X sky130_fd_sc_hd__mux2_1
XFILLER_138_1305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12347_ _17889_/Q _12347_/B vssd1 vssd1 vccd1 vccd1 _12348_/A sky130_fd_sc_hd__and2_1
XFILLER_114_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15066_ _15083_/A vssd1 vssd1 vccd1 vccd1 _15066_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_142_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12278_ _11530_/A _11512_/C _17874_/Q vssd1 vssd1 vccd1 vccd1 _12279_/B sky130_fd_sc_hd__o21bai_1
X_14017_ _14017_/A vssd1 vssd1 vccd1 vccd1 _14017_/X sky130_fd_sc_hd__buf_6
XFILLER_4_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11229_ _11232_/A _11232_/C vssd1 vssd1 vccd1 vccd1 _11231_/A sky130_fd_sc_hd__and2_1
XFILLER_96_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_214_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18825_ _18860_/CLK _18825_/D vssd1 vssd1 vccd1 vccd1 _18825_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_68_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18756_ _18786_/CLK _18756_/D vssd1 vssd1 vccd1 vccd1 _18756_/Q sky130_fd_sc_hd__dfxtp_2
X_15968_ _16000_/A _15971_/B vssd1 vssd1 vccd1 vccd1 _15968_/Y sky130_fd_sc_hd__nand2_1
XTAP_5490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17707_ _09509_/Y _13356_/B _13363_/Y _18990_/Q vssd1 vssd1 vccd1 vccd1 _18990_/D
+ sky130_fd_sc_hd__a22o_1
X_14919_ _14919_/A _15371_/B _14965_/C vssd1 vssd1 vccd1 vccd1 _14919_/X sky130_fd_sc_hd__or3_1
XFILLER_110_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18687_ _18693_/CLK _18687_/D vssd1 vssd1 vccd1 vccd1 _18687_/Q sky130_fd_sc_hd__dfxtp_2
X_15899_ _18590_/Q _18554_/Q _15899_/S vssd1 vssd1 vccd1 vccd1 _15899_/X sky130_fd_sc_hd__mux2_1
XFILLER_58_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_1366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_224_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17638_ _17638_/A _17638_/B vssd1 vssd1 vccd1 vccd1 _17639_/A sky130_fd_sc_hd__and2_1
XFILLER_145_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_184_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17569_ _17587_/A _17569_/B vssd1 vssd1 vccd1 vccd1 _17570_/A sky130_fd_sc_hd__and2_1
XFILLER_210_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_204_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_177_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_192_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_1260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09825_ _17782_/Q vssd1 vssd1 vccd1 vccd1 _11032_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_86_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09756_ _18096_/Q _17978_/Q vssd1 vssd1 vccd1 vccd1 _10611_/B sky130_fd_sc_hd__xor2_4
XFILLER_230_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_189_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09687_ _10575_/B vssd1 vssd1 vccd1 vccd1 _09688_/A sky130_fd_sc_hd__buf_6
XTAP_2116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_214_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10600_ _10600_/A _10600_/B vssd1 vssd1 vccd1 vccd1 _10600_/X sky130_fd_sc_hd__or2_1
XFILLER_167_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11580_ _11842_/A _11502_/X _11537_/Y _11579_/X vssd1 vssd1 vccd1 vccd1 _11680_/A
+ sky130_fd_sc_hd__o31a_1
XFILLER_10_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10531_ _10529_/X _10530_/X _10926_/A vssd1 vssd1 vccd1 vccd1 _10531_/X sky130_fd_sc_hd__mux2_2
XFILLER_10_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13250_ _13250_/A vssd1 vssd1 vccd1 vccd1 _18078_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_6_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10462_ _10521_/A vssd1 vssd1 vccd1 vccd1 _10462_/X sky130_fd_sc_hd__buf_6
XFILLER_182_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_202_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12201_ _17853_/Q _11709_/B _17854_/Q vssd1 vssd1 vccd1 vccd1 _12201_/X sky130_fd_sc_hd__a21o_1
X_13181_ _13181_/A vssd1 vssd1 vccd1 vccd1 _18047_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_108_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10393_ _10333_/S _10390_/X _10392_/X _09965_/A vssd1 vssd1 vccd1 vccd1 _10393_/X
+ sky130_fd_sc_hd__o31a_1
XFILLER_191_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12132_ _12132_/A _12132_/B _12132_/C _12132_/D vssd1 vssd1 vccd1 vccd1 _12132_/X
+ sky130_fd_sc_hd__or4_2
XFILLER_123_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16940_ _16999_/A vssd1 vssd1 vccd1 vccd1 _16940_/X sky130_fd_sc_hd__clkbuf_2
X_12063_ _12063_/A _12102_/B vssd1 vssd1 vccd1 vccd1 _12069_/B sky130_fd_sc_hd__xnor2_1
XFILLER_150_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11014_ _17996_/Q vssd1 vssd1 vccd1 vccd1 _13375_/C sky130_fd_sc_hd__buf_2
XFILLER_89_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_1295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16871_ _16871_/A vssd1 vssd1 vccd1 vccd1 _16871_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_131_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18610_ _18614_/CLK _18610_/D vssd1 vssd1 vccd1 vccd1 _18610_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_37_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15822_ _15857_/A _16128_/B _15870_/C vssd1 vssd1 vccd1 vccd1 _15822_/X sky130_fd_sc_hd__or3_1
XTAP_4030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_213_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_219_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18541_ _18542_/CLK _18541_/D vssd1 vssd1 vccd1 vccd1 _18541_/Q sky130_fd_sc_hd__dfxtp_2
X_15753_ _18554_/Q _18518_/Q _15753_/S vssd1 vssd1 vccd1 vccd1 _15753_/X sky130_fd_sc_hd__mux2_1
XTAP_4074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_218_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_80 _13591_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12965_ _12958_/A _12952_/X _12963_/X _12964_/X vssd1 vssd1 vccd1 vccd1 _17974_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_64_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINSDIODE2_91 _13752_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14704_ _18178_/Q _18177_/Q _14704_/C vssd1 vssd1 vccd1 vccd1 _15145_/C sky130_fd_sc_hd__or3_4
X_11916_ _11916_/A _11916_/B vssd1 vssd1 vccd1 vccd1 _11917_/B sky130_fd_sc_hd__nor2_1
X_15684_ _18500_/Q _15683_/B _15683_/Y _15681_/X vssd1 vssd1 vccd1 vccd1 _18500_/D
+ sky130_fd_sc_hd__o211a_1
X_18472_ _18473_/CLK _18472_/D vssd1 vssd1 vccd1 vccd1 _18472_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_3384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12896_ _17960_/Q _12792_/X _12890_/B _17962_/Q vssd1 vssd1 vccd1 vccd1 _12897_/C
+ sky130_fd_sc_hd__a31o_1
XTAP_2650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_206_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14635_ _14683_/A _14635_/B vssd1 vssd1 vccd1 vccd1 _14635_/Y sky130_fd_sc_hd__nand2_1
XFILLER_54_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17423_ _17423_/A _17538_/C vssd1 vssd1 vccd1 vccd1 _17432_/B sky130_fd_sc_hd__nor2_2
X_11847_ _11621_/Y _11846_/X _11635_/X vssd1 vssd1 vccd1 vccd1 _11850_/C sky130_fd_sc_hd__a21oi_1
XTAP_2694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_221_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_159_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14566_ _16835_/A vssd1 vssd1 vccd1 vccd1 _15172_/A sky130_fd_sc_hd__buf_8
XTAP_1993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17354_ _17376_/A _17493_/B _17376_/C vssd1 vssd1 vccd1 vccd1 _17354_/X sky130_fd_sc_hd__or3_1
X_11778_ _11774_/Y _11777_/X _11781_/A _11776_/Y vssd1 vssd1 vccd1 vccd1 _11778_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_41_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16305_ _16329_/A _16305_/B vssd1 vssd1 vccd1 vccd1 _16305_/Y sky130_fd_sc_hd__nand2_1
X_13517_ _18675_/Q _13493_/X _13500_/X _18690_/Q _13516_/X vssd1 vssd1 vccd1 vccd1
+ _13517_/X sky130_fd_sc_hd__a221o_1
XFILLER_53_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10729_ _09109_/A _10737_/S _10728_/X _10743_/A vssd1 vssd1 vccd1 vccd1 _10729_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_146_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17285_ _18919_/Q _18883_/Q _17298_/S vssd1 vssd1 vccd1 vccd1 _17285_/X sky130_fd_sc_hd__mux2_1
X_14497_ _14497_/A vssd1 vssd1 vccd1 vccd1 _18222_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_173_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_174_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_220_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16236_ _18666_/Q _18630_/Q _16250_/S vssd1 vssd1 vccd1 vccd1 _16236_/X sky130_fd_sc_hd__mux2_1
XFILLER_118_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19024_ _19026_/CLK _19024_/D vssd1 vssd1 vccd1 vccd1 _19024_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_70_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13448_ _13448_/A vssd1 vssd1 vccd1 vccd1 _13448_/Y sky130_fd_sc_hd__inv_2
XFILLER_9_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_220_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16167_ _16922_/A vssd1 vssd1 vccd1 vccd1 _16759_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_173_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13379_ _17768_/A _13379_/B _13379_/C vssd1 vssd1 vccd1 vccd1 _13380_/A sky130_fd_sc_hd__and3_1
XFILLER_127_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15118_ _15118_/A _15118_/B vssd1 vssd1 vccd1 vccd1 _15118_/Y sky130_fd_sc_hd__nand2_1
Xclkbuf_4_7_0_wb_clk_i clkbuf_4_7_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_4_7_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_5_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16098_ _16096_/B _16095_/X _16096_/Y _16097_/X vssd1 vssd1 vccd1 vccd1 _18599_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_126_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_1321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15049_ _15061_/A _15049_/B vssd1 vssd1 vccd1 vccd1 _15049_/Y sky130_fd_sc_hd__nand2_1
XFILLER_214_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_229_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_229_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_214_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_44_wb_clk_i clkbuf_5_16_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18812_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_96_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09610_ _09610_/A _09610_/B vssd1 vssd1 vccd1 vccd1 _09611_/B sky130_fd_sc_hd__xnor2_4
X_18808_ _18809_/CLK _18808_/D vssd1 vssd1 vccd1 vccd1 _18808_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_56_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_209_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09541_ _09589_/B _09541_/B vssd1 vssd1 vccd1 vccd1 _10007_/B sky130_fd_sc_hd__or2_2
X_18739_ _18743_/CLK _18739_/D vssd1 vssd1 vccd1 vccd1 _18739_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_37_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09472_ _09472_/A vssd1 vssd1 vccd1 vccd1 _18142_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_37_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_221_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_221_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_211_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_221_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_146_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_145_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_219_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09808_ _09808_/A _09808_/B vssd1 vssd1 vccd1 vccd1 _09810_/A sky130_fd_sc_hd__xnor2_1
XFILLER_87_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09739_ _09739_/A _09739_/B vssd1 vssd1 vccd1 vccd1 _09752_/B sky130_fd_sc_hd__xnor2_1
XFILLER_189_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12750_ _18029_/Q _18028_/Q _18031_/Q _18030_/Q vssd1 vssd1 vccd1 vccd1 _12752_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_216_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11701_ _11701_/A vssd1 vssd1 vccd1 vccd1 _11848_/A sky130_fd_sc_hd__clkbuf_2
XTAP_1234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_215_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_187_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12681_ _12676_/B _12613_/A _12679_/Y _12680_/X _12667_/X vssd1 vssd1 vccd1 vccd1
+ _17933_/D sky130_fd_sc_hd__a221o_1
XTAP_1256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14420_ _14420_/A _14420_/B vssd1 vssd1 vccd1 vccd1 _18195_/D sky130_fd_sc_hd__nor2_1
XTAP_1289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11632_ _11681_/D _11730_/B vssd1 vssd1 vccd1 vccd1 _11633_/B sky130_fd_sc_hd__nand2_1
XFILLER_42_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_230_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14351_ _18995_/Q _10982_/X _14272_/X _14350_/X vssd1 vssd1 vccd1 vccd1 _18181_/D
+ sky130_fd_sc_hd__o2bb2a_1
X_11563_ _19032_/Q _11563_/B _11563_/C vssd1 vssd1 vccd1 vccd1 _11563_/X sky130_fd_sc_hd__and3_1
XFILLER_156_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13302_ _18050_/Q _18053_/Q _18052_/Q _18055_/Q vssd1 vssd1 vccd1 vccd1 _13303_/C
+ sky130_fd_sc_hd__or4_1
XFILLER_195_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17070_ _17503_/A _17070_/B vssd1 vssd1 vccd1 vccd1 _17080_/B sky130_fd_sc_hd__nor2_2
X_10514_ _11925_/A _10506_/X _10510_/X _10512_/X _10903_/S vssd1 vssd1 vccd1 vccd1
+ _10515_/C sky130_fd_sc_hd__a311o_1
XFILLER_13_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14282_ _14282_/A vssd1 vssd1 vccd1 vccd1 _14282_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_11494_ _11654_/B _11788_/A vssd1 vssd1 vccd1 vccd1 _13444_/A sky130_fd_sc_hd__nor2_1
XFILLER_109_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16021_ _16043_/A _16021_/B _16021_/C vssd1 vssd1 vccd1 vccd1 _16021_/X sky130_fd_sc_hd__or3_1
XFILLER_137_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13233_ _13233_/A _18072_/Q vssd1 vssd1 vccd1 vccd1 _13234_/A sky130_fd_sc_hd__and2_1
XFILLER_7_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10445_ _09248_/C _09253_/D _10503_/S vssd1 vssd1 vccd1 vccd1 _10445_/X sky130_fd_sc_hd__mux2_1
XFILLER_170_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13164_ _13164_/A _18041_/Q vssd1 vssd1 vccd1 vccd1 _13165_/A sky130_fd_sc_hd__and2_1
XFILLER_156_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10376_ _10782_/A _10376_/B vssd1 vssd1 vccd1 vccd1 _10376_/X sky130_fd_sc_hd__or2_1
XFILLER_83_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_124_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12115_ _10829_/X _09828_/B _12114_/X vssd1 vssd1 vccd1 vccd1 _12116_/B sky130_fd_sc_hd__a21o_1
XFILLER_97_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13095_ _17709_/A _18008_/Q vssd1 vssd1 vccd1 vccd1 _13096_/A sky130_fd_sc_hd__or2_1
X_17972_ _18108_/CLK _17972_/D vssd1 vssd1 vccd1 vccd1 _17972_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_215_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16923_ _16936_/A _17506_/B _16936_/C vssd1 vssd1 vccd1 vccd1 _16923_/X sky130_fd_sc_hd__or3_1
XFILLER_133_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12046_ _12047_/A _12133_/B vssd1 vssd1 vccd1 vccd1 _12054_/A sky130_fd_sc_hd__and2_1
XFILLER_133_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16854_ _16866_/A _17449_/B _16866_/C vssd1 vssd1 vccd1 vccd1 _16854_/X sky130_fd_sc_hd__or3_1
XFILLER_92_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15805_ _18566_/Q _18530_/Q _15809_/S vssd1 vssd1 vccd1 vccd1 _15805_/X sky130_fd_sc_hd__mux2_1
XFILLER_225_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13997_ _18586_/Q _13738_/A _13995_/X _13996_/X vssd1 vssd1 vccd1 vccd1 _13997_/X
+ sky130_fd_sc_hd__a211o_1
X_16785_ _16796_/A _16785_/B _16796_/C vssd1 vssd1 vccd1 vccd1 _16785_/X sky130_fd_sc_hd__or3_1
XFILLER_46_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18524_ _18532_/CLK _18524_/D vssd1 vssd1 vccd1 vccd1 _18524_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_18_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15736_ _15736_/A vssd1 vssd1 vccd1 vccd1 _15753_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_19_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12948_ _18036_/Q _13310_/A _12948_/C vssd1 vssd1 vccd1 vccd1 _12948_/X sky130_fd_sc_hd__and3_1
XFILLER_74_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_206_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_162_wb_clk_i _18114_/CLK vssd1 vssd1 vccd1 vccd1 _18108_/CLK sky130_fd_sc_hd__clkbuf_16
X_18455_ _18458_/CLK _18455_/D vssd1 vssd1 vccd1 vccd1 _18455_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_209_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15667_ _15673_/B _15665_/X _15666_/X _15662_/X vssd1 vssd1 vccd1 vccd1 _18495_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_179_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12879_ _12881_/B _12888_/B _12879_/C vssd1 vssd1 vccd1 vccd1 _12880_/A sky130_fd_sc_hd__and3b_1
XTAP_2480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_222_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17406_ _18950_/Q _18914_/Q _17406_/S vssd1 vssd1 vccd1 vccd1 _17406_/X sky130_fd_sc_hd__mux2_1
XFILLER_178_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14618_ _17556_/A vssd1 vssd1 vccd1 vccd1 _14618_/X sky130_fd_sc_hd__buf_2
X_18386_ _18387_/CLK _18386_/D vssd1 vssd1 vccd1 vccd1 _18386_/Q sky130_fd_sc_hd__dfxtp_4
X_15598_ _18516_/Q _18480_/Q _15604_/S vssd1 vssd1 vccd1 vccd1 _15598_/X sky130_fd_sc_hd__mux2_1
XFILLER_92_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14549_ _14637_/A vssd1 vssd1 vccd1 vccd1 _17635_/A sky130_fd_sc_hd__clkbuf_2
X_17337_ _18896_/Q _17336_/B _17336_/Y _17324_/X vssd1 vssd1 vccd1 vccd1 _18896_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_202_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_222_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17268_ _17448_/A vssd1 vssd1 vccd1 vccd1 _17318_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_101_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19007_ _19009_/CLK _19007_/D vssd1 vssd1 vccd1 vccd1 _19007_/Q sky130_fd_sc_hd__dfxtp_1
X_16219_ _16219_/A vssd1 vssd1 vccd1 vccd1 _16807_/A sky130_fd_sc_hd__buf_6
XFILLER_161_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_220_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17199_ _18899_/Q _18863_/Q _17199_/S vssd1 vssd1 vccd1 vccd1 _17199_/X sky130_fd_sc_hd__mux2_1
XFILLER_115_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_103_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08972_ _08972_/A vssd1 vssd1 vccd1 vccd1 _08972_/Y sky130_fd_sc_hd__inv_2
XFILLER_216_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_1260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_216_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_217_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09524_ _18992_/Q vssd1 vssd1 vccd1 vccd1 _14199_/A sky130_fd_sc_hd__inv_2
XFILLER_71_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_231_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_227_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_213_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09455_ _09272_/A _09440_/Y _09466_/B vssd1 vssd1 vccd1 vccd1 _09475_/B sky130_fd_sc_hd__a21o_1
XPHY_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_227_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_212_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_185_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09386_ _09386_/A _09386_/B _09972_/A _09386_/D vssd1 vssd1 vccd1 vccd1 _09387_/C
+ sky130_fd_sc_hd__and4_1
XFILLER_200_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_1294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_197_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_180_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_193_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10230_ _10518_/A vssd1 vssd1 vccd1 vccd1 _10489_/S sky130_fd_sc_hd__buf_2
XFILLER_3_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10161_ _10141_/A _10141_/B _10160_/X vssd1 vssd1 vccd1 vccd1 _10168_/B sky130_fd_sc_hd__o21bai_2
XFILLER_126_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10092_ _10086_/Y _10091_/Y _12061_/A vssd1 vssd1 vccd1 vccd1 _10092_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13920_ _18754_/Q _14124_/A _13706_/X _18736_/Q vssd1 vssd1 vccd1 vccd1 _13920_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_130_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13851_ _18703_/Q _13591_/X _13592_/X _18727_/Q vssd1 vssd1 vccd1 vccd1 _13851_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_19_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12802_ _17956_/Q vssd1 vssd1 vccd1 vccd1 _12802_/Y sky130_fd_sc_hd__inv_2
XFILLER_90_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13782_ _18432_/Q _13847_/A _13781_/X _18423_/Q vssd1 vssd1 vccd1 vccd1 _13782_/X
+ sky130_fd_sc_hd__a22o_1
X_16570_ _16621_/A vssd1 vssd1 vccd1 vccd1 _16598_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_74_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_222_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10994_ _17778_/Q _09518_/B _09517_/Y vssd1 vssd1 vccd1 vccd1 _17778_/D sky130_fd_sc_hd__a21o_1
XFILLER_90_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15521_ _15566_/A _15525_/B vssd1 vssd1 vccd1 vccd1 _15521_/Y sky130_fd_sc_hd__nand2_1
XFILLER_128_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12733_ _19024_/Q _19023_/Q _19026_/Q _19025_/Q vssd1 vssd1 vccd1 vccd1 _12736_/A
+ sky130_fd_sc_hd__and4_1
XTAP_1031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_206_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_187_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_231_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_204_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15452_ _15516_/A vssd1 vssd1 vccd1 vccd1 _15452_/X sky130_fd_sc_hd__clkbuf_2
X_18240_ _18245_/CLK _18240_/D vssd1 vssd1 vccd1 vccd1 _18240_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12664_ _12656_/A _12656_/B _12654_/A vssd1 vssd1 vccd1 vccd1 _12665_/B sky130_fd_sc_hd__a21o_1
XFILLER_230_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_1178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_141_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14403_ _14420_/A _14403_/B vssd1 vssd1 vccd1 vccd1 _18191_/D sky130_fd_sc_hd__nor2_1
XFILLER_175_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11615_ _11615_/A _17858_/Q vssd1 vssd1 vccd1 vccd1 _11615_/Y sky130_fd_sc_hd__nor2_1
X_15383_ _15390_/B _15379_/X _15381_/X _15382_/X vssd1 vssd1 vccd1 vccd1 _18429_/D
+ sky130_fd_sc_hd__o211a_1
X_18171_ _18184_/CLK _18171_/D vssd1 vssd1 vccd1 vccd1 _18171_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12595_ _17924_/Q vssd1 vssd1 vccd1 vccd1 _12597_/B sky130_fd_sc_hd__clkinv_2
XFILLER_129_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_184_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17122_ _17412_/A _17256_/C vssd1 vssd1 vccd1 vccd1 _17129_/B sky130_fd_sc_hd__nor2_2
X_14334_ _14334_/A _14334_/B vssd1 vssd1 vccd1 vccd1 _14334_/Y sky130_fd_sc_hd__nor2_1
XFILLER_129_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11546_ _11546_/A _11546_/B _11546_/C vssd1 vssd1 vccd1 vccd1 _11621_/B sky130_fd_sc_hd__and3_1
XFILLER_102_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17053_ _17088_/A _17056_/B vssd1 vssd1 vccd1 vccd1 _17053_/Y sky130_fd_sc_hd__nand2_1
X_14265_ _10985_/X _12085_/B _14237_/X _12097_/B vssd1 vssd1 vccd1 vccd1 _14265_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_167_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11477_ _11459_/A _12337_/S _11338_/A _11479_/B vssd1 vssd1 vccd1 vccd1 _11477_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_137_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16004_ _16003_/B _16002_/X _16003_/Y _15988_/X vssd1 vssd1 vccd1 vccd1 _18578_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_125_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13216_ _13222_/A _18064_/Q vssd1 vssd1 vccd1 vccd1 _13217_/A sky130_fd_sc_hd__and2_1
XFILLER_109_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10428_ _10560_/S vssd1 vssd1 vccd1 vccd1 _10494_/A sky130_fd_sc_hd__buf_2
XFILLER_143_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14196_ _14196_/A _14196_/B _14196_/C vssd1 vssd1 vccd1 vccd1 _14216_/B sky130_fd_sc_hd__or3_2
XFILLER_140_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13147_ _13151_/A _18033_/Q vssd1 vssd1 vccd1 vccd1 _13148_/A sky130_fd_sc_hd__and2_1
XTAP_815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10359_ _10366_/B _10403_/A vssd1 vssd1 vccd1 vccd1 _10605_/C sky130_fd_sc_hd__and2_1
XTAP_826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13078_ _13076_/X _13077_/X _12346_/A vssd1 vssd1 vccd1 vccd1 _13078_/Y sky130_fd_sc_hd__a21oi_1
X_17955_ _17959_/CLK _17955_/D vssd1 vssd1 vccd1 vccd1 _17955_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_97_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16906_ _17491_/A _16906_/B vssd1 vssd1 vccd1 vccd1 _16916_/B sky130_fd_sc_hd__nor2_2
X_12029_ _12055_/D _12029_/B vssd1 vssd1 vccd1 vccd1 _12099_/B sky130_fd_sc_hd__or2_4
X_17886_ _17890_/CLK _17886_/D vssd1 vssd1 vccd1 vccd1 _17886_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_18_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_226_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16837_ _17435_/A _16906_/B vssd1 vssd1 vccd1 vccd1 _16847_/B sky130_fd_sc_hd__nor2_2
XFILLER_38_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16768_ _16832_/A vssd1 vssd1 vccd1 vccd1 _16815_/A sky130_fd_sc_hd__clkbuf_2
X_18507_ _18511_/CLK _18507_/D vssd1 vssd1 vccd1 vccd1 _18507_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_34_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_206_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15719_ _15754_/A _15719_/B vssd1 vssd1 vccd1 vccd1 _15719_/Y sky130_fd_sc_hd__nand2_1
XFILLER_20_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16699_ _16699_/A _16699_/B vssd1 vssd1 vccd1 vccd1 _16699_/Y sky130_fd_sc_hd__nand2_1
XFILLER_55_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_222_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_146_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09240_ _18905_/Q _18904_/Q _18903_/Q vssd1 vssd1 vccd1 vccd1 _09243_/B sky130_fd_sc_hd__or3_4
X_18438_ _18443_/CLK _18438_/D vssd1 vssd1 vccd1 vccd1 _18438_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_146_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_222_1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09171_ _09171_/A _09171_/B _09171_/C vssd1 vssd1 vccd1 vccd1 _09188_/A sky130_fd_sc_hd__and3_1
X_18369_ _18374_/CLK _18369_/D vssd1 vssd1 vccd1 vccd1 _18369_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_175_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_159_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_5_16_0_wb_clk_i clkbuf_4_8_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_5_16_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_143_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08955_ _08967_/A vssd1 vssd1 vccd1 vccd1 _08960_/A sky130_fd_sc_hd__buf_12
XTAP_5319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_116_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_217_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_217_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_204_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09507_ _17591_/A _14383_/B vssd1 vssd1 vccd1 vccd1 _17704_/A sky130_fd_sc_hd__nand2_1
XFILLER_225_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_198_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_213_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_197_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09438_ _09475_/A _09467_/A vssd1 vssd1 vccd1 vccd1 _09439_/A sky130_fd_sc_hd__or2_1
XFILLER_52_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_212_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_169_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09369_ _18281_/Q _18280_/Q _18279_/Q vssd1 vssd1 vccd1 vccd1 _10883_/A sky130_fd_sc_hd__or3_2
XFILLER_205_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11400_ _11466_/B _11467_/C _11307_/B _11467_/D vssd1 vssd1 vccd1 vccd1 _11442_/B
+ sky130_fd_sc_hd__a31o_1
X_12380_ _12380_/A vssd1 vssd1 vccd1 vccd1 _17894_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_122_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11331_ _17878_/Q _19030_/Q vssd1 vssd1 vccd1 vccd1 _11331_/X sky130_fd_sc_hd__or2b_1
XFILLER_107_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_197_1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14050_ _12055_/A _14042_/X _14049_/X _13684_/Y vssd1 vssd1 vccd1 vccd1 _14050_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_158_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11262_ _17800_/Q _11287_/A _11261_/X vssd1 vssd1 vccd1 vccd1 _12036_/B sky130_fd_sc_hd__a21o_1
XFILLER_107_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_106_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13001_ _13001_/A _13005_/B vssd1 vssd1 vccd1 vccd1 _13001_/Y sky130_fd_sc_hd__nor2_1
XFILLER_107_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10213_ _10213_/A _10213_/B vssd1 vssd1 vccd1 vccd1 _10218_/B sky130_fd_sc_hd__xnor2_1
XFILLER_133_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_1305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11193_ _11196_/B _11193_/B vssd1 vssd1 vccd1 vccd1 _11194_/B sky130_fd_sc_hd__xnor2_1
XFILLER_84_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10144_ _10144_/A _10148_/B vssd1 vssd1 vccd1 vccd1 _10146_/B sky130_fd_sc_hd__xor2_1
XFILLER_122_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17740_ _17740_/A vssd1 vssd1 vccd1 vccd1 _19013_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14952_ _18363_/Q _18327_/Q _14955_/S vssd1 vssd1 vccd1 vccd1 _14952_/X sky130_fd_sc_hd__mux2_1
X_10075_ _09103_/A _09098_/D _09093_/D _09103_/C _09995_/A _09708_/A vssd1 vssd1 vccd1
+ vccd1 _10075_/X sky130_fd_sc_hd__mux4_1
XFILLER_94_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13903_ _18538_/Q _13705_/A _13902_/X vssd1 vssd1 vccd1 vccd1 _13903_/X sky130_fd_sc_hd__a21o_1
XFILLER_48_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17671_ _17645_/X _17663_/Y _17654_/X _17664_/Y _18980_/Q vssd1 vssd1 vccd1 vccd1
+ _17672_/B sky130_fd_sc_hd__a32o_1
X_14883_ _18346_/Q _18310_/Q _14883_/S vssd1 vssd1 vccd1 vccd1 _14883_/X sky130_fd_sc_hd__mux2_1
XFILLER_90_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16622_ _18761_/Q _18725_/Q _16637_/S vssd1 vssd1 vccd1 vccd1 _16622_/X sky130_fd_sc_hd__mux2_1
XFILLER_35_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13834_ _13834_/A vssd1 vssd1 vccd1 vccd1 _13834_/X sky130_fd_sc_hd__buf_6
XINSDIODE2_205 _13066_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_223_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XINSDIODE2_216 _13723_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_216_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XINSDIODE2_227 _15175_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16553_ _16701_/A _16602_/B vssd1 vssd1 vccd1 vccd1 _16562_/B sky130_fd_sc_hd__nor2_1
XINSDIODE2_238 _18413_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13765_ _18486_/Q _13735_/X _13764_/X _18510_/Q vssd1 vssd1 vccd1 vccd1 _13765_/X
+ sky130_fd_sc_hd__a22o_1
XPHY_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XINSDIODE2_249 _09098_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10977_ _10977_/A vssd1 vssd1 vccd1 vccd1 _10977_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_31_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15504_ _15562_/A vssd1 vssd1 vccd1 vccd1 _15551_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_188_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_206_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_204_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12716_ _13019_/B vssd1 vssd1 vccd1 vccd1 _12951_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_203_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16484_ _16507_/A _16487_/B vssd1 vssd1 vccd1 vccd1 _16484_/Y sky130_fd_sc_hd__nand2_1
XFILLER_15_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13696_ _13649_/X _13662_/X _13695_/X _14507_/B vssd1 vssd1 vccd1 vccd1 _13696_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_231_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18223_ _19026_/CLK _18223_/D vssd1 vssd1 vccd1 vccd1 _18223_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_15_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15435_ _18477_/Q _18441_/Q _15435_/S vssd1 vssd1 vccd1 vccd1 _15435_/X sky130_fd_sc_hd__mux2_1
XFILLER_175_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12647_ _12647_/A _12647_/B vssd1 vssd1 vccd1 vccd1 _12649_/A sky130_fd_sc_hd__nor2_1
XFILLER_19_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15366_ _15375_/A _15366_/B vssd1 vssd1 vccd1 vccd1 _15366_/Y sky130_fd_sc_hd__nand2_1
XFILLER_175_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18154_ _18157_/CLK _18154_/D vssd1 vssd1 vccd1 vccd1 _18154_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_7_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12578_ _17921_/Q _12569_/X _12576_/X _12577_/Y _12548_/X vssd1 vssd1 vccd1 vccd1
+ _17921_/D sky130_fd_sc_hd__a221o_1
XFILLER_172_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17105_ _17156_/A _17105_/B vssd1 vssd1 vccd1 vccd1 _17105_/Y sky130_fd_sc_hd__nand2_1
XFILLER_171_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11529_ _17873_/Q vssd1 vssd1 vccd1 vccd1 _11530_/A sky130_fd_sc_hd__inv_2
X_14317_ _14317_/A _14317_/B vssd1 vssd1 vccd1 vccd1 _14317_/Y sky130_fd_sc_hd__nand2_1
X_15297_ _15370_/A vssd1 vssd1 vccd1 vccd1 _15448_/B sky130_fd_sc_hd__buf_2
XFILLER_184_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_183_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18085_ _18085_/CLK _18085_/D vssd1 vssd1 vccd1 vccd1 _18085_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_7_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17036_ _17035_/B _17034_/X _17035_/Y _17020_/X vssd1 vssd1 vccd1 vccd1 _18821_/D
+ sky130_fd_sc_hd__o211a_1
X_14248_ _10985_/X _09657_/X _14205_/X _11924_/A _14247_/Y vssd1 vssd1 vccd1 vccd1
+ _14248_/X sky130_fd_sc_hd__a221o_1
XFILLER_132_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_217_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14179_ _18668_/Q _13508_/X _14177_/X _14178_/X vssd1 vssd1 vccd1 vccd1 _14179_/X
+ sky130_fd_sc_hd__a211o_1
XTAP_601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18987_ _18989_/CLK _18987_/D vssd1 vssd1 vccd1 vccd1 _18987_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_227_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17938_ _17939_/CLK _17938_/D vssd1 vssd1 vccd1 vccd1 _17938_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_26_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_226_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_187_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_1293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_227_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17869_ _19032_/CLK _17869_/D vssd1 vssd1 vccd1 vccd1 _17869_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_94_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_226_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_187_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_226_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_228_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_224_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09223_ _18947_/Q _18946_/Q _18945_/Q vssd1 vssd1 vccd1 vccd1 _09227_/A sky130_fd_sc_hd__or3_4
XFILLER_195_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09154_ _09154_/A _09154_/B _09154_/C vssd1 vssd1 vccd1 vccd1 _09429_/A sky130_fd_sc_hd__and3_1
XFILLER_33_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09085_ _17838_/Q _17837_/Q _17835_/Q vssd1 vssd1 vccd1 vccd1 _09086_/A sky130_fd_sc_hd__and3_4
X_19116__87 vssd1 vssd1 vccd1 vccd1 _19116__87/HI _19224_/A sky130_fd_sc_hd__conb_1
XFILLER_162_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_104_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09987_ _09987_/A vssd1 vssd1 vccd1 vccd1 _09987_/X sky130_fd_sc_hd__buf_4
XTAP_5127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08938_ _08941_/A vssd1 vssd1 vccd1 vccd1 _08938_/Y sky130_fd_sc_hd__inv_2
XTAP_5149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10900_ _09413_/A _09408_/C _09418_/D _10956_/A _10542_/X _10518_/X vssd1 vssd1 vccd1
+ vccd1 _10900_/X sky130_fd_sc_hd__mux4_2
XFILLER_85_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11880_ _13094_/A vssd1 vssd1 vccd1 vccd1 _13210_/A sky130_fd_sc_hd__buf_4
XTAP_3769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10831_ _10829_/X _10830_/X _10689_/A vssd1 vssd1 vccd1 vccd1 _10831_/X sky130_fd_sc_hd__a21o_1
XFILLER_16_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13550_ _13940_/A vssd1 vssd1 vccd1 vccd1 _13837_/A sky130_fd_sc_hd__buf_6
XFILLER_13_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10762_ _09186_/C _09176_/B _10883_/B vssd1 vssd1 vccd1 vccd1 _10762_/X sky130_fd_sc_hd__mux2_1
XFILLER_16_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_213_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12501_ _17910_/Q _12492_/A _12484_/X _12500_/X vssd1 vssd1 vccd1 vccd1 _12501_/X
+ sky130_fd_sc_hd__o31a_1
XFILLER_12_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13481_ _14421_/A vssd1 vssd1 vccd1 vccd1 _14420_/A sky130_fd_sc_hd__buf_4
XFILLER_51_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10693_ _10811_/A vssd1 vssd1 vccd1 vccd1 _10693_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_13_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15220_ _15220_/A _15220_/B _15257_/C vssd1 vssd1 vccd1 vccd1 _15220_/X sky130_fd_sc_hd__or3_1
XFILLER_12_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12432_ _12459_/A _12432_/B _12432_/C vssd1 vssd1 vccd1 vccd1 _12433_/A sky130_fd_sc_hd__and3_1
XFILLER_201_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15151_ _18375_/Q _15154_/B _15150_/X _15143_/X vssd1 vssd1 vccd1 vccd1 _18375_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_138_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12363_ _12467_/C vssd1 vssd1 vccd1 vccd1 _12472_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_201_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14102_ _18635_/Q _14017_/A _14098_/X _14101_/X vssd1 vssd1 vccd1 vccd1 _14102_/X
+ sky130_fd_sc_hd__a211o_1
X_11314_ _11337_/A _11313_/X _11297_/Y vssd1 vssd1 vccd1 vccd1 _11375_/B sky130_fd_sc_hd__a21boi_1
X_15082_ _15118_/A _15082_/B vssd1 vssd1 vccd1 vccd1 _15082_/Y sky130_fd_sc_hd__nand2_1
XFILLER_180_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12294_ _12294_/A vssd1 vssd1 vccd1 vccd1 _17872_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_49_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14033_ _18263_/Q _13838_/A _14031_/X _14032_/X vssd1 vssd1 vccd1 vccd1 _14033_/X
+ sky130_fd_sc_hd__a211o_1
X_18910_ _18927_/CLK _18910_/D vssd1 vssd1 vccd1 vccd1 _18910_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_153_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11245_ _11245_/A _11245_/B vssd1 vssd1 vccd1 vccd1 _11245_/Y sky130_fd_sc_hd__nand2_1
XFILLER_171_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_1274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18841_ _18845_/CLK _18841_/D vssd1 vssd1 vccd1 vccd1 _18841_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_164_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11176_ _17806_/Q _17805_/Q _11212_/B vssd1 vssd1 vccd1 vccd1 _11184_/C sky130_fd_sc_hd__and3_1
XFILLER_110_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10127_ _10181_/A vssd1 vssd1 vccd1 vccd1 _10440_/A sky130_fd_sc_hd__clkinv_4
X_18772_ _18773_/CLK _18772_/D vssd1 vssd1 vccd1 vccd1 _18772_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_95_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15984_ _15984_/A _15984_/B _16021_/C vssd1 vssd1 vccd1 vccd1 _15984_/X sky130_fd_sc_hd__or3_1
XTAP_5661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17723_ _17723_/A _19007_/Q vssd1 vssd1 vccd1 vccd1 _17724_/A sky130_fd_sc_hd__and2_1
XTAP_5683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14935_ _14935_/A _14935_/B vssd1 vssd1 vccd1 vccd1 _14935_/Y sky130_fd_sc_hd__nand2_1
X_10058_ _10010_/A _10054_/X _10057_/X vssd1 vssd1 vccd1 vccd1 _10058_/X sky130_fd_sc_hd__a21o_1
XFILLER_57_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_224_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17654_ _17675_/A vssd1 vssd1 vccd1 vccd1 _17654_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_4993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14866_ _14958_/A vssd1 vssd1 vccd1 vccd1 _14883_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_35_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16605_ _16615_/A _16749_/B _16628_/C vssd1 vssd1 vccd1 vccd1 _16605_/X sky130_fd_sc_hd__or3_1
XFILLER_17_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_223_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13817_ _18933_/Q _13785_/X _13815_/X _13816_/X vssd1 vssd1 vccd1 vccd1 _13817_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_17_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17585_ _17585_/A vssd1 vssd1 vccd1 vccd1 _18958_/D sky130_fd_sc_hd__clkbuf_1
X_14797_ _15840_/A vssd1 vssd1 vccd1 vccd1 _15207_/A sky130_fd_sc_hd__buf_2
XFILLER_51_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_1340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_69_wb_clk_i clkbuf_opt_1_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18732_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_16_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16536_ _16538_/B _16534_/X _16535_/Y _16519_/X vssd1 vssd1 vccd1 vccd1 _18703_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_204_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13748_ _13434_/A _13729_/X _13747_/X _12055_/A vssd1 vssd1 vccd1 vccd1 _13829_/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_16_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_177_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16467_ _18723_/Q _18687_/Q _16470_/S vssd1 vssd1 vccd1 vccd1 _16467_/X sky130_fd_sc_hd__mux2_1
XFILLER_177_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13679_ _18522_/Q _13677_/X _13623_/A _18528_/Q _13678_/X vssd1 vssd1 vccd1 vccd1
+ _13679_/X sky130_fd_sc_hd__a221o_1
XFILLER_85_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18206_ _18992_/CLK _18206_/D vssd1 vssd1 vccd1 vccd1 _18206_/Q sky130_fd_sc_hd__dfxtp_1
X_15418_ _15417_/B _15416_/X _15417_/Y _15404_/X vssd1 vssd1 vccd1 vccd1 _18437_/D
+ sky130_fd_sc_hd__o211a_1
X_19186_ _19186_/A _09002_/Y vssd1 vssd1 vccd1 vccd1 io_out[24] sky130_fd_sc_hd__ebufn_8
X_16398_ _16456_/A vssd1 vssd1 vccd1 vccd1 _16398_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_185_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18137_ _18140_/CLK _18137_/D vssd1 vssd1 vccd1 vccd1 _18137_/Q sky130_fd_sc_hd__dfxtp_1
X_15349_ _15373_/A _15352_/B vssd1 vssd1 vccd1 vccd1 _15349_/Y sky130_fd_sc_hd__nand2_1
XFILLER_172_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18068_ _18068_/CLK _18068_/D vssd1 vssd1 vccd1 vccd1 _18068_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_208_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17019_ _17323_/A vssd1 vssd1 vccd1 vccd1 _17096_/A sky130_fd_sc_hd__clkbuf_2
X_09910_ _09902_/A _09910_/B vssd1 vssd1 vccd1 vccd1 _09962_/A sky130_fd_sc_hd__and2b_1
XFILLER_217_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09841_ _09855_/A _09855_/B _09840_/X vssd1 vssd1 vccd1 vccd1 _09842_/B sky130_fd_sc_hd__o21ba_1
XFILLER_113_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_217_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_1366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09772_ _09781_/A _09781_/B vssd1 vssd1 vccd1 vccd1 _09774_/B sky130_fd_sc_hd__xnor2_4
XFILLER_218_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_224_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_226_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_214_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_226_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09206_ _18680_/Q _18679_/Q _18678_/Q vssd1 vssd1 vccd1 vccd1 _09209_/B sky130_fd_sc_hd__or3_4
XFILLER_139_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09137_ _09137_/A _09137_/B _09137_/C vssd1 vssd1 vccd1 vccd1 _09138_/B sky130_fd_sc_hd__and3_1
XFILLER_147_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_159_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09068_ _09068_/A vssd1 vssd1 vccd1 vccd1 _19177_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_191_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11030_ _17972_/Q _11036_/B vssd1 vssd1 vccd1 vccd1 _13337_/A sky130_fd_sc_hd__or2_1
XFILLER_104_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12981_ _12967_/A _12958_/B _12980_/X vssd1 vssd1 vccd1 vccd1 _12982_/B sky130_fd_sc_hd__a21oi_1
XFILLER_64_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14720_ _14833_/A vssd1 vssd1 vccd1 vccd1 _14812_/A sky130_fd_sc_hd__buf_2
XTAP_3533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11932_ _11932_/A _11976_/A vssd1 vssd1 vccd1 vccd1 _11983_/A sky130_fd_sc_hd__nand2_1
XTAP_3555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_5_9_0_wb_clk_i clkbuf_5_9_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_5_9_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_72_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14651_ _14651_/A _15241_/A vssd1 vssd1 vccd1 vccd1 _14658_/B sky130_fd_sc_hd__nor2_1
XTAP_3588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11863_ _17764_/A vssd1 vssd1 vccd1 vccd1 _11863_/X sky130_fd_sc_hd__buf_4
XTAP_3599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13602_ _18732_/Q _13575_/X _13576_/X _18723_/Q _13601_/X vssd1 vssd1 vccd1 vccd1
+ _13602_/X sky130_fd_sc_hd__a221o_2
X_10814_ _09270_/A _10687_/A _10813_/X _10770_/X vssd1 vssd1 vccd1 vccd1 _10814_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_2887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_220_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17370_ _17370_/A vssd1 vssd1 vccd1 vccd1 _17386_/S sky130_fd_sc_hd__clkbuf_2
XTAP_2898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14582_ _16850_/A vssd1 vssd1 vccd1 vccd1 _16853_/A sky130_fd_sc_hd__buf_8
X_11794_ _11749_/B _11786_/Y _11787_/X _11729_/X _11793_/X vssd1 vssd1 vccd1 vccd1
+ _11794_/X sky130_fd_sc_hd__o221a_1
XFILLER_186_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16321_ _16503_/A vssd1 vssd1 vccd1 vccd1 _16371_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_13533_ _13552_/B _13541_/B vssd1 vssd1 vccd1 vccd1 _13724_/A sky130_fd_sc_hd__nor2_1
X_10745_ _09114_/C _10350_/A _10841_/A vssd1 vssd1 vccd1 vccd1 _10745_/X sky130_fd_sc_hd__mux2_1
XFILLER_129_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_199_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16252_ _16252_/A vssd1 vssd1 vccd1 vccd1 _16252_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_13464_ _13456_/B _13455_/A _13457_/A vssd1 vssd1 vccd1 vccd1 _13464_/X sky130_fd_sc_hd__a21o_1
XFILLER_139_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10676_ _12102_/A _12101_/A vssd1 vssd1 vccd1 vccd1 _10833_/A sky130_fd_sc_hd__and2_1
XFILLER_90_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15203_ _15236_/A _15206_/B vssd1 vssd1 vccd1 vccd1 _15203_/Y sky130_fd_sc_hd__nand2_1
X_12415_ _12413_/X _12415_/B _12467_/C vssd1 vssd1 vccd1 vccd1 _12416_/A sky130_fd_sc_hd__and3b_1
XFILLER_51_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16183_ _18655_/Q _18619_/Q _16192_/S vssd1 vssd1 vccd1 vccd1 _16183_/X sky130_fd_sc_hd__mux2_1
X_13395_ _13405_/B vssd1 vssd1 vccd1 vccd1 _13395_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_86_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15134_ _15277_/A _15134_/B vssd1 vssd1 vccd1 vccd1 _15142_/B sky130_fd_sc_hd__nor2_2
X_12346_ _12346_/A _12346_/B _12346_/C vssd1 vssd1 vccd1 vccd1 _17888_/D sky130_fd_sc_hd__nor3_1
XFILLER_182_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_187_wb_clk_i clkbuf_5_8_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17884_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_5_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_116_wb_clk_i clkbuf_5_30_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18469_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_15065_ _15098_/A _15371_/B _15112_/C vssd1 vssd1 vccd1 vccd1 _15065_/X sky130_fd_sc_hd__or3_1
X_12277_ _12277_/A vssd1 vssd1 vccd1 vccd1 _17869_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_218_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14016_ _14016_/A vssd1 vssd1 vccd1 vccd1 _14017_/A sky130_fd_sc_hd__buf_6
X_11228_ _11228_/A vssd1 vssd1 vccd1 vccd1 _17818_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_214_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18824_ _18858_/CLK _18824_/D vssd1 vssd1 vccd1 vccd1 _18824_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_68_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11159_ _11780_/A _17814_/Q _12285_/A vssd1 vssd1 vccd1 vccd1 _11160_/A sky130_fd_sc_hd__mux2_1
XFILLER_68_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18755_ _18788_/CLK _18755_/D vssd1 vssd1 vccd1 vccd1 _18755_/Q sky130_fd_sc_hd__dfxtp_2
X_15967_ _18604_/Q _18568_/Q _15990_/S vssd1 vssd1 vccd1 vccd1 _15967_/X sky130_fd_sc_hd__mux2_1
XTAP_5480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17706_ _17706_/A vssd1 vssd1 vccd1 vccd1 _18989_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_208_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14918_ _14918_/A vssd1 vssd1 vccd1 vccd1 _14965_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_3_1349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18686_ _18686_/CLK _18686_/D vssd1 vssd1 vccd1 vccd1 _18686_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_82_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15898_ _15900_/B _15896_/X _15897_/Y _15881_/X vssd1 vssd1 vccd1 vccd1 _18553_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_4790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17637_ _17575_/X _17635_/Y _17631_/X _17636_/Y _18972_/Q vssd1 vssd1 vccd1 vccd1
+ _17638_/B sky130_fd_sc_hd__a32o_1
X_14849_ _14875_/A _14849_/B vssd1 vssd1 vccd1 vccd1 _14849_/Y sky130_fd_sc_hd__nand2_1
XFILLER_1_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_225_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_223_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17568_ _17567_/X _17560_/Y _17561_/X _17562_/Y _18955_/Q vssd1 vssd1 vccd1 vccd1
+ _17569_/B sky130_fd_sc_hd__a32o_1
XFILLER_51_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_225_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16519_ _16559_/A vssd1 vssd1 vccd1 vccd1 _16519_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_20_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_220_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17499_ _17519_/A vssd1 vssd1 vccd1 vccd1 _17515_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_143_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_219_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19169_ _19169_/A _09016_/Y vssd1 vssd1 vccd1 vccd1 io_out[7] sky130_fd_sc_hd__ebufn_8
XFILLER_118_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_1272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09824_ _09843_/A _12112_/A vssd1 vssd1 vccd1 vccd1 _09855_/A sky130_fd_sc_hd__nand2_2
XFILLER_98_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09755_ _18102_/Q _10116_/B vssd1 vssd1 vccd1 vccd1 _09760_/A sky130_fd_sc_hd__xnor2_2
XFILLER_228_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09686_ _09991_/A vssd1 vssd1 vccd1 vccd1 _10575_/B sky130_fd_sc_hd__buf_2
XTAP_2106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_227_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_230_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_214_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_202_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_211_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_196_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10530_ _09165_/A _09160_/C _09170_/D _10308_/A _10484_/A _10489_/S vssd1 vssd1 vccd1
+ vccd1 _10530_/X sky130_fd_sc_hd__mux4_1
XFILLER_183_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_155_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10461_ _11924_/A _10453_/X _10460_/X _12039_/A vssd1 vssd1 vccd1 vccd1 _10461_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_148_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12200_ _12205_/A vssd1 vssd1 vccd1 vccd1 _12200_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_108_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13180_ _13186_/A _18048_/Q vssd1 vssd1 vccd1 vccd1 _13181_/A sky130_fd_sc_hd__and2_1
XFILLER_202_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_202_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10392_ _09344_/B _09950_/X _10391_/X _09969_/A vssd1 vssd1 vccd1 vccd1 _10392_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_163_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12131_ _12131_/A _13635_/A vssd1 vssd1 vccd1 vccd1 _12132_/D sky130_fd_sc_hd__xor2_1
XFILLER_11_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12062_ _10948_/S _12092_/B _12060_/X _12061_/X vssd1 vssd1 vccd1 vccd1 _12069_/A
+ sky130_fd_sc_hd__a211o_1
XFILLER_111_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_0_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_1_0_1_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_132_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11013_ _17997_/Q vssd1 vssd1 vccd1 vccd1 _13375_/B sky130_fd_sc_hd__buf_2
XFILLER_132_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16870_ _16882_/A _16874_/B vssd1 vssd1 vccd1 vccd1 _16870_/Y sky130_fd_sc_hd__nand2_1
XFILLER_49_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19100__71 vssd1 vssd1 vccd1 vccd1 _19100__71/HI _19208_/A sky130_fd_sc_hd__conb_1
XFILLER_78_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15821_ _15821_/A vssd1 vssd1 vccd1 vccd1 _15870_/C sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_4020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18540_ _18542_/CLK _18540_/D vssd1 vssd1 vccd1 vccd1 _18540_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_4064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15752_ _15754_/B _15750_/X _15751_/Y _15740_/X vssd1 vssd1 vccd1 vccd1 _18517_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_4075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_70 _13523_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12964_ _13037_/A vssd1 vssd1 vccd1 vccd1 _12964_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_79_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XINSDIODE2_81 _13591_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_92 _13670_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14703_ _16219_/A vssd1 vssd1 vccd1 vccd1 _15292_/A sky130_fd_sc_hd__buf_4
XTAP_3363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18471_ _18473_/CLK _18471_/D vssd1 vssd1 vccd1 vccd1 _18471_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_3374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11915_ _12982_/A _11915_/B vssd1 vssd1 vccd1 vccd1 _11918_/A sky130_fd_sc_hd__xnor2_1
X_15683_ _15694_/A _15683_/B vssd1 vssd1 vccd1 vccd1 _15683_/Y sky130_fd_sc_hd__nand2_1
XFILLER_206_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12895_ _17961_/Q _17962_/Q _12895_/C vssd1 vssd1 vccd1 vccd1 _12899_/B sky130_fd_sc_hd__and3_1
XTAP_2651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17422_ _18917_/Q _17419_/B _17419_/Y _17421_/X vssd1 vssd1 vccd1 vccd1 _18917_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_205_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14634_ _17544_/A vssd1 vssd1 vccd1 vccd1 _14683_/A sky130_fd_sc_hd__buf_2
XTAP_2673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11846_ _11609_/X _11617_/X _11848_/A vssd1 vssd1 vccd1 vccd1 _11846_/X sky130_fd_sc_hd__a21o_1
XTAP_2684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_159_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_1204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17353_ _18936_/Q _18900_/Q _17367_/S vssd1 vssd1 vccd1 vccd1 _17353_/X sky130_fd_sc_hd__mux2_1
X_11777_ _11781_/A _11776_/Y _11769_/X _11772_/X vssd1 vssd1 vccd1 vccd1 _11777_/X
+ sky130_fd_sc_hd__o2bb2a_1
X_14565_ _14593_/A _17674_/A vssd1 vssd1 vccd1 vccd1 _16835_/A sky130_fd_sc_hd__or2_4
XFILLER_14_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16304_ _18683_/Q _18647_/Q _16304_/S vssd1 vssd1 vccd1 vccd1 _16304_/X sky130_fd_sc_hd__mux2_1
X_13516_ _18666_/Q _13508_/X _13515_/X _18672_/Q vssd1 vssd1 vccd1 vccd1 _13516_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_147_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10728_ _10728_/A _10763_/S vssd1 vssd1 vccd1 vccd1 _10728_/X sky130_fd_sc_hd__or2_1
X_17284_ _17291_/B _17281_/X _17282_/X _17283_/X vssd1 vssd1 vccd1 vccd1 _18882_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_140_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14496_ _18222_/Q _14502_/B vssd1 vssd1 vccd1 vccd1 _14497_/A sky130_fd_sc_hd__and2_1
XFILLER_146_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19023_ _19026_/CLK _19023_/D vssd1 vssd1 vccd1 vccd1 _19023_/Q sky130_fd_sc_hd__dfxtp_1
X_16235_ _16327_/A vssd1 vssd1 vccd1 vccd1 _16250_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_220_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10659_ _10812_/S vssd1 vssd1 vccd1 vccd1 _10858_/S sky130_fd_sc_hd__buf_4
XFILLER_139_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13447_ _13447_/A _13447_/B vssd1 vssd1 vccd1 vccd1 _13447_/X sky130_fd_sc_hd__or2_1
XFILLER_155_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_220_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16166_ _18651_/Q _18615_/Q _16170_/S vssd1 vssd1 vccd1 vccd1 _16166_/X sky130_fd_sc_hd__mux2_1
X_13378_ _10113_/A _13337_/A _13368_/Y vssd1 vssd1 vccd1 vccd1 _13379_/C sky130_fd_sc_hd__a21o_1
XFILLER_142_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15117_ _18404_/Q _18368_/Q _15121_/S vssd1 vssd1 vccd1 vccd1 _15117_/X sky130_fd_sc_hd__mux2_1
XFILLER_170_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12329_ _12329_/A _12329_/B _12329_/C vssd1 vssd1 vccd1 vccd1 _12330_/C sky130_fd_sc_hd__nand3_1
X_16097_ _16139_/A vssd1 vssd1 vccd1 vccd1 _16097_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_173_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15048_ _18386_/Q _18350_/Q _15052_/S vssd1 vssd1 vccd1 vccd1 _15048_/X sky130_fd_sc_hd__mux2_1
XFILLER_190_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_1355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_229_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_205_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_1358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18807_ _18809_/CLK _18807_/D vssd1 vssd1 vccd1 vccd1 _18807_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_28_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16999_ _16999_/A vssd1 vssd1 vccd1 vccd1 _16999_/X sky130_fd_sc_hd__clkbuf_2
Xclkbuf_leaf_84_wb_clk_i _18144_/CLK vssd1 vssd1 vccd1 vccd1 _18620_/CLK sky130_fd_sc_hd__clkbuf_16
X_09540_ _10181_/A _09540_/B vssd1 vssd1 vccd1 vccd1 _09541_/B sky130_fd_sc_hd__nor2_1
X_18738_ _18738_/CLK _18738_/D vssd1 vssd1 vccd1 vccd1 _18738_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_23_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_224_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_13_wb_clk_i clkbuf_5_4_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17969_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_09471_ _09482_/A _09471_/B vssd1 vssd1 vccd1 vccd1 _09472_/A sky130_fd_sc_hd__or2_1
XFILLER_58_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18669_ _18686_/CLK _18669_/D vssd1 vssd1 vccd1 vccd1 _18669_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_52_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_97_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_149_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_211_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_225_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_221_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_165_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_166_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_161_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_219_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09807_ _09807_/A _09807_/B vssd1 vssd1 vccd1 vccd1 _09808_/B sky130_fd_sc_hd__xnor2_1
XFILLER_132_1280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09738_ _18111_/Q vssd1 vssd1 vccd1 vccd1 _09752_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_28_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_227_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09669_ _09639_/B _09669_/B vssd1 vssd1 vccd1 vccd1 _09669_/X sky130_fd_sc_hd__and2b_1
XFILLER_83_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_231_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11700_ _11700_/A _11706_/A vssd1 vssd1 vccd1 vccd1 _11700_/Y sky130_fd_sc_hd__nor2_1
XTAP_1224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12680_ _12679_/A _12679_/B _12537_/S vssd1 vssd1 vccd1 vccd1 _12680_/X sky130_fd_sc_hd__o21a_1
XFILLER_76_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11631_ _11621_/Y _11627_/Y _11630_/X _11390_/X vssd1 vssd1 vccd1 vccd1 _11631_/X
+ sky130_fd_sc_hd__o22a_1
XTAP_1268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_91_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_168_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11562_ _11562_/A _17866_/Q vssd1 vssd1 vccd1 vccd1 _11563_/C sky130_fd_sc_hd__nor2_1
X_14350_ _15607_/C _14349_/Y _17709_/A vssd1 vssd1 vccd1 vccd1 _14350_/X sky130_fd_sc_hd__a21o_1
XFILLER_128_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_204_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13301_ _18038_/Q _18041_/Q _18040_/Q _18043_/Q vssd1 vssd1 vccd1 vccd1 _13303_/B
+ sky130_fd_sc_hd__or4_1
XFILLER_10_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10513_ _10513_/A vssd1 vssd1 vccd1 vccd1 _10903_/S sky130_fd_sc_hd__buf_2
X_14281_ _14203_/X _14293_/A _14296_/A _14280_/Y vssd1 vssd1 vccd1 vccd1 _14281_/X
+ sky130_fd_sc_hd__o22a_1
X_11493_ _11446_/X _11451_/Y _11492_/X vssd1 vssd1 vccd1 vccd1 _11493_/X sky130_fd_sc_hd__a21o_1
XFILLER_155_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16020_ _18618_/Q _18582_/Q _16031_/S vssd1 vssd1 vccd1 vccd1 _16020_/X sky130_fd_sc_hd__mux2_1
XFILLER_171_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13232_ _13232_/A vssd1 vssd1 vccd1 vccd1 _18070_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_109_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10444_ _10494_/A vssd1 vssd1 vccd1 vccd1 _10503_/S sky130_fd_sc_hd__buf_4
XFILLER_137_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13163_ _13163_/A vssd1 vssd1 vccd1 vccd1 _18039_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_48_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10375_ _09332_/A _09337_/B _10375_/S vssd1 vssd1 vccd1 vccd1 _10375_/X sky130_fd_sc_hd__mux2_1
XFILLER_3_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_152_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12114_ _10829_/X _09828_/B _11032_/A vssd1 vssd1 vccd1 vccd1 _12114_/X sky130_fd_sc_hd__o21a_1
XFILLER_135_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13094_ _13094_/A vssd1 vssd1 vccd1 vccd1 _17709_/A sky130_fd_sc_hd__buf_4
X_17971_ _18108_/CLK _17971_/D vssd1 vssd1 vccd1 vccd1 _17971_/Q sky130_fd_sc_hd__dfxtp_1
X_19077__48 vssd1 vssd1 vccd1 vccd1 _19077__48/HI _19171_/A sky130_fd_sc_hd__conb_1
XFILLER_46_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16922_ _16922_/A vssd1 vssd1 vccd1 vccd1 _17506_/B sky130_fd_sc_hd__buf_6
X_12045_ _12101_/B vssd1 vssd1 vccd1 vccd1 _12133_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_105_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_172_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16853_ _16853_/A vssd1 vssd1 vccd1 vccd1 _17449_/B sky130_fd_sc_hd__buf_4
XFILLER_172_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15804_ _15806_/B _15801_/X _15802_/Y _15803_/X vssd1 vssd1 vccd1 vccd1 _18529_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_168_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16784_ _18801_/Q _18765_/Q _16784_/S vssd1 vssd1 vccd1 vccd1 _16784_/X sky130_fd_sc_hd__mux2_1
XFILLER_219_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13996_ _18574_/Q _13785_/A _13743_/A _18556_/Q vssd1 vssd1 vccd1 vccd1 _13996_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_19_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18523_ _18532_/CLK _18523_/D vssd1 vssd1 vccd1 vccd1 _18523_/Q sky130_fd_sc_hd__dfxtp_4
X_15735_ _15743_/B _15733_/X _15734_/X _15720_/X vssd1 vssd1 vccd1 vccd1 _18513_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_20_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12947_ _12947_/A _12983_/A vssd1 vssd1 vccd1 vccd1 _12947_/X sky130_fd_sc_hd__or2_1
XFILLER_65_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18454_ _18458_/CLK _18454_/D vssd1 vssd1 vccd1 vccd1 _18454_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_222_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15666_ _15678_/A _15964_/B _15666_/C vssd1 vssd1 vccd1 vccd1 _15666_/X sky130_fd_sc_hd__or3_1
XFILLER_61_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12878_ _17954_/Q _12824_/A _12869_/A _17956_/Q vssd1 vssd1 vccd1 vccd1 _12879_/C
+ sky130_fd_sc_hd__a31o_1
XTAP_2481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17405_ _17408_/B _17402_/X _17404_/Y _17400_/X vssd1 vssd1 vccd1 vccd1 _18913_/D
+ sky130_fd_sc_hd__o211a_1
X_14617_ _14584_/B _14612_/A _18248_/Q vssd1 vssd1 vccd1 vccd1 _14617_/Y sky130_fd_sc_hd__o21bai_1
X_18385_ _18387_/CLK _18385_/D vssd1 vssd1 vccd1 vccd1 _18385_/Q sky130_fd_sc_hd__dfxtp_4
X_11829_ _11705_/D _11714_/B _11828_/Y vssd1 vssd1 vccd1 vccd1 _11829_/X sky130_fd_sc_hd__o21a_1
XFILLER_60_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15597_ _16041_/A _15597_/B vssd1 vssd1 vccd1 vccd1 _15605_/B sky130_fd_sc_hd__nor2_2
XFILLER_21_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_222_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_221_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_202_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17336_ _17336_/A _17336_/B vssd1 vssd1 vccd1 vccd1 _17336_/Y sky130_fd_sc_hd__nand2_1
XFILLER_186_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14548_ _18174_/Q _18173_/Q _18170_/Q _18169_/Q vssd1 vssd1 vccd1 vccd1 _14637_/A
+ sky130_fd_sc_hd__or4b_2
XFILLER_147_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_131_wb_clk_i clkbuf_5_24_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18406_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_186_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17267_ _17412_/A _17399_/C vssd1 vssd1 vccd1 vccd1 _17275_/B sky130_fd_sc_hd__nor2_2
XFILLER_140_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14479_ _14479_/A vssd1 vssd1 vccd1 vccd1 _18214_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_31_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19006_ _19009_/CLK _19006_/D vssd1 vssd1 vccd1 vccd1 _19006_/Q sky130_fd_sc_hd__dfxtp_1
X_16218_ _16217_/B _16215_/X _16217_/Y _16209_/X vssd1 vssd1 vccd1 vccd1 _18626_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_220_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17198_ _17200_/B _17195_/X _17196_/Y _17197_/X vssd1 vssd1 vccd1 vccd1 _18862_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_128_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16149_ _16905_/A vssd1 vssd1 vccd1 vccd1 _16745_/A sky130_fd_sc_hd__buf_6
XFILLER_143_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08971_ _08972_/A vssd1 vssd1 vccd1 vccd1 _08971_/Y sky130_fd_sc_hd__inv_2
XFILLER_216_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_1272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_229_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_69_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19091__62 vssd1 vssd1 vccd1 vccd1 _19091__62/HI _19199_/A sky130_fd_sc_hd__conb_1
XFILLER_83_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09523_ _10990_/A vssd1 vssd1 vccd1 vccd1 _09523_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_71_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_225_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_224_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_225_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09454_ _09138_/B _09454_/B _09454_/C vssd1 vssd1 vccd1 vccd1 _09466_/B sky130_fd_sc_hd__and3b_1
XFILLER_149_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09385_ _18404_/Q _18403_/Q _18402_/Q vssd1 vssd1 vccd1 vccd1 _09386_/D sky130_fd_sc_hd__or3_4
Xclkbuf_leaf_219_wb_clk_i _17864_/CLK vssd1 vssd1 vccd1 vccd1 _19032_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_101_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_184_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_220_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_203_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_158_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10160_ _10140_/A _10160_/B vssd1 vssd1 vccd1 vccd1 _10160_/X sky130_fd_sc_hd__and2b_1
XFILLER_160_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10091_ _10044_/A _10087_/X _10090_/X _10009_/A vssd1 vssd1 vccd1 vccd1 _10091_/Y
+ sky130_fd_sc_hd__a22oi_2
XFILLER_82_1274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13850_ _18715_/Q _13581_/X _13582_/X _18709_/Q _13849_/X vssd1 vssd1 vccd1 vccd1
+ _13850_/X sky130_fd_sc_hd__a221o_1
XFILLER_142_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12801_ _17916_/Q _12839_/A _12798_/Y _17937_/Q _12800_/X vssd1 vssd1 vccd1 vccd1
+ _12813_/A sky130_fd_sc_hd__a221o_1
XFILLER_142_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_210_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13781_ _13781_/A vssd1 vssd1 vccd1 vccd1 _13781_/X sky130_fd_sc_hd__clkbuf_16
X_10993_ _17778_/Q _09509_/Y _09518_/X _17780_/Q vssd1 vssd1 vccd1 vccd1 _17780_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_27_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15520_ _15578_/A vssd1 vssd1 vccd1 vccd1 _15566_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_204_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12732_ _12987_/A _13310_/A vssd1 vssd1 vccd1 vccd1 _13318_/C sky130_fd_sc_hd__and2_1
XFILLER_76_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_231_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15451_ _15492_/A _16043_/B _15451_/C vssd1 vssd1 vccd1 vccd1 _15451_/X sky130_fd_sc_hd__or3_1
XFILLER_187_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12663_ _12663_/A _12663_/B vssd1 vssd1 vccd1 vccd1 _12665_/A sky130_fd_sc_hd__nor2_1
XFILLER_203_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14402_ _18191_/Q _14398_/Y _14401_/X _09495_/B vssd1 vssd1 vccd1 vccd1 _14403_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_187_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11614_ _11614_/A _12221_/A vssd1 vssd1 vccd1 vccd1 _11614_/Y sky130_fd_sc_hd__nand2_1
XFILLER_30_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18170_ _18184_/CLK _18170_/D vssd1 vssd1 vccd1 vccd1 _18170_/Q sky130_fd_sc_hd__dfxtp_1
X_15382_ _15404_/A vssd1 vssd1 vccd1 vccd1 _15382_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_141_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12594_ _12629_/A _12594_/B vssd1 vssd1 vccd1 vccd1 _12600_/A sky130_fd_sc_hd__nand2_1
XFILLER_211_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_196_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17121_ _17184_/A vssd1 vssd1 vccd1 vccd1 _17256_/C sky130_fd_sc_hd__buf_2
XFILLER_184_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14333_ _14334_/A _14334_/B vssd1 vssd1 vccd1 vccd1 _14333_/X sky130_fd_sc_hd__and2_1
X_11545_ _11617_/A _11617_/B _12089_/B vssd1 vssd1 vccd1 vccd1 _11546_/C sky130_fd_sc_hd__o21ai_1
X_17052_ _18862_/Q _18826_/Q _17055_/S vssd1 vssd1 vccd1 vccd1 _17052_/X sky130_fd_sc_hd__mux2_1
XFILLER_13_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11476_ _11525_/B _11474_/X _11475_/X vssd1 vssd1 vccd1 vccd1 _11476_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_7_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14264_ _14202_/X _14262_/X _14263_/X _13334_/X vssd1 vssd1 vccd1 vccd1 _18172_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_100_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16003_ _16003_/A _16003_/B vssd1 vssd1 vccd1 vccd1 _16003_/Y sky130_fd_sc_hd__nand2_1
XFILLER_100_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13215_ _13215_/A vssd1 vssd1 vccd1 vccd1 _18062_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_48_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10427_ _10899_/A _10427_/B vssd1 vssd1 vccd1 vccd1 _10427_/X sky130_fd_sc_hd__and2_1
XFILLER_171_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14195_ _18214_/Q _18213_/Q _18212_/Q vssd1 vssd1 vccd1 vccd1 _14196_/C sky130_fd_sc_hd__or3_2
XFILLER_125_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10358_ _10346_/X _10353_/X _10357_/X _09981_/X vssd1 vssd1 vccd1 vccd1 _10358_/X
+ sky130_fd_sc_hd__o31a_1
X_13146_ _13146_/A vssd1 vssd1 vccd1 vccd1 _18031_/D sky130_fd_sc_hd__clkbuf_1
XTAP_805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13077_ _18005_/Q _18006_/Q vssd1 vssd1 vccd1 vccd1 _13077_/X sky130_fd_sc_hd__xor2_1
X_17954_ _17954_/CLK _17954_/D vssd1 vssd1 vccd1 vccd1 _17954_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_61_1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_183_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10289_ _09969_/X _10281_/Y _10288_/Y _12128_/A vssd1 vssd1 vccd1 vccd1 _10289_/Y
+ sky130_fd_sc_hd__a211oi_2
X_12028_ _12028_/A _12028_/B _12028_/C _12028_/D vssd1 vssd1 vccd1 vccd1 _12029_/B
+ sky130_fd_sc_hd__or4_1
X_16905_ _16905_/A vssd1 vssd1 vccd1 vccd1 _17491_/A sky130_fd_sc_hd__buf_4
XFILLER_111_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17885_ _17888_/CLK _17885_/D vssd1 vssd1 vccd1 vccd1 _17885_/Q sky130_fd_sc_hd__dfxtp_1
X_16836_ _16879_/A vssd1 vssd1 vccd1 vccd1 _16906_/B sky130_fd_sc_hd__buf_2
XFILLER_65_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16767_ _18797_/Q _18761_/Q _16784_/S vssd1 vssd1 vccd1 vccd1 _16767_/X sky130_fd_sc_hd__mux2_1
XFILLER_4_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13979_ _18361_/Q _13559_/A _13772_/X _18355_/Q _13978_/X vssd1 vssd1 vccd1 vccd1
+ _13979_/X sky130_fd_sc_hd__a221o_1
XFILLER_34_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_206_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18506_ _18506_/CLK _18506_/D vssd1 vssd1 vccd1 vccd1 _18506_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_207_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15718_ _18545_/Q _18509_/Q _15733_/S vssd1 vssd1 vccd1 vccd1 _15718_/X sky130_fd_sc_hd__mux2_1
XFILLER_20_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16698_ _18779_/Q _18743_/Q _16715_/S vssd1 vssd1 vccd1 vccd1 _16698_/X sky130_fd_sc_hd__mux2_1
XFILLER_94_1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18437_ _18443_/CLK _18437_/D vssd1 vssd1 vccd1 vccd1 _18437_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_34_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15649_ _15649_/A vssd1 vssd1 vccd1 vccd1 _15889_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_94_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_178_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_203_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09170_ _09170_/A _09170_/B _09170_/C _09170_/D vssd1 vssd1 vccd1 vccd1 _09171_/C
+ sky130_fd_sc_hd__and4_1
XFILLER_21_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18368_ _18380_/CLK _18368_/D vssd1 vssd1 vccd1 vccd1 _18368_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_222_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17319_ _17327_/B _17317_/X _17318_/X _17304_/X vssd1 vssd1 vccd1 vccd1 _18891_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_119_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_186_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18299_ _18299_/CLK _18299_/D vssd1 vssd1 vccd1 vccd1 _18299_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_175_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_190_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_128_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08954_ _08954_/A vssd1 vssd1 vccd1 vccd1 _08954_/Y sky130_fd_sc_hd__inv_2
XFILLER_69_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_217_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_227_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09506_ _18205_/Q _09506_/B vssd1 vssd1 vccd1 vccd1 _14383_/B sky130_fd_sc_hd__or2_2
XFILLER_25_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_227_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_212_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09437_ _09482_/A _09474_/A vssd1 vssd1 vccd1 vccd1 _09467_/A sky130_fd_sc_hd__or2_1
XFILLER_53_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09368_ _18296_/Q _18295_/Q _18294_/Q vssd1 vssd1 vccd1 vccd1 _09370_/C sky130_fd_sc_hd__or3_4
XFILLER_40_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_197_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09299_ _10569_/A _09299_/B _09299_/C _09299_/D vssd1 vssd1 vccd1 vccd1 _09299_/X
+ sky130_fd_sc_hd__and4_1
XFILLER_201_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_177_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11330_ _11345_/A vssd1 vssd1 vccd1 vccd1 _11330_/Y sky130_fd_sc_hd__inv_2
XFILLER_193_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_193_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11261_ _17802_/Q _17801_/Q vssd1 vssd1 vccd1 vccd1 _11261_/X sky130_fd_sc_hd__or2_2
XFILLER_197_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13000_ _13000_/A _13000_/B _13000_/C vssd1 vssd1 vccd1 vccd1 _13005_/B sky130_fd_sc_hd__and3_1
X_10212_ _13372_/A vssd1 vssd1 vccd1 vccd1 _10218_/A sky130_fd_sc_hd__inv_2
XFILLER_107_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11192_ _11192_/A vssd1 vssd1 vccd1 vccd1 _17809_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_171_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_1328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10143_ _18127_/Q _10118_/B _10142_/Y vssd1 vssd1 vccd1 vccd1 _10148_/B sky130_fd_sc_hd__a21o_1
X_19047__18 vssd1 vssd1 vccd1 vccd1 _19047__18/HI _19141_/A sky130_fd_sc_hd__conb_1
XTAP_5810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14951_ _15241_/A _14985_/B vssd1 vssd1 vccd1 vccd1 _14960_/B sky130_fd_sc_hd__nor2_2
X_10074_ _09098_/A _09093_/C _09103_/D _09098_/B _09987_/A _09708_/A vssd1 vssd1 vccd1
+ vccd1 _10074_/X sky130_fd_sc_hd__mux4_1
XFILLER_94_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13902_ _18523_/Q _13505_/A _13734_/A _18529_/Q vssd1 vssd1 vccd1 vccd1 _13902_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_5887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17670_ _17670_/A vssd1 vssd1 vccd1 vccd1 _18979_/D sky130_fd_sc_hd__clkbuf_1
XTAP_5898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14882_ _14890_/B _14879_/X _14880_/X _14881_/X vssd1 vssd1 vccd1 vccd1 _18309_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_169_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16621_ _16621_/A vssd1 vssd1 vccd1 vccd1 _16637_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_47_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13833_ _13833_/A vssd1 vssd1 vccd1 vccd1 _18166_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_90_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_206 _12862_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XINSDIODE2_217 _13730_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16552_ _16551_/B _16550_/X _16551_/Y _16539_/X vssd1 vssd1 vccd1 vccd1 _18707_/D
+ sky130_fd_sc_hd__o211a_1
X_13764_ _13764_/A vssd1 vssd1 vccd1 vccd1 _13764_/X sky130_fd_sc_hd__clkbuf_4
XINSDIODE2_228 _15199_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_239 _18358_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10976_ _14222_/A _14272_/B vssd1 vssd1 vccd1 vccd1 _10977_/A sky130_fd_sc_hd__nand2_1
X_15503_ _18492_/Q _18456_/Q _15514_/S vssd1 vssd1 vccd1 vccd1 _15503_/X sky130_fd_sc_hd__mux2_1
X_12715_ _12748_/A vssd1 vssd1 vccd1 vccd1 _13019_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_71_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_188_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16483_ _18727_/Q _18691_/Q _16490_/S vssd1 vssd1 vccd1 vccd1 _16483_/X sky130_fd_sc_hd__mux2_1
X_13695_ _12027_/A _13675_/X _13683_/X _13684_/Y _13694_/X vssd1 vssd1 vccd1 vccd1
+ _13695_/X sky130_fd_sc_hd__a221o_1
XFILLER_204_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18222_ _18222_/CLK _18222_/D vssd1 vssd1 vccd1 vccd1 _18222_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_231_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15434_ _16030_/A _15448_/B vssd1 vssd1 vccd1 vccd1 _15445_/B sky130_fd_sc_hd__nor2_2
XFILLER_148_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12646_ _12646_/A _12646_/B vssd1 vssd1 vccd1 vccd1 _12647_/B sky130_fd_sc_hd__nor2_1
XFILLER_203_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_157_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18153_ _19000_/CLK _18153_/D vssd1 vssd1 vccd1 vccd1 _18153_/Q sky130_fd_sc_hd__dfxtp_1
X_15365_ _18461_/Q _18425_/Q _15388_/S vssd1 vssd1 vccd1 vccd1 _15365_/X sky130_fd_sc_hd__mux2_1
XFILLER_184_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12577_ _12561_/Y _12575_/Y _12571_/X _12569_/A vssd1 vssd1 vccd1 vccd1 _12577_/Y
+ sky130_fd_sc_hd__a31oi_1
XFILLER_50_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17104_ _17168_/A vssd1 vssd1 vccd1 vccd1 _17156_/A sky130_fd_sc_hd__buf_2
XFILLER_7_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14316_ _14275_/X _14313_/X _14315_/X _14270_/X vssd1 vssd1 vccd1 vccd1 _18177_/D
+ sky130_fd_sc_hd__o211a_1
X_11528_ _11732_/A _11528_/B _11410_/A vssd1 vssd1 vccd1 vccd1 _11528_/X sky130_fd_sc_hd__or3b_1
X_18084_ _18087_/CLK _18084_/D vssd1 vssd1 vccd1 vccd1 _18084_/Q sky130_fd_sc_hd__dfxtp_1
X_15296_ _16219_/A vssd1 vssd1 vccd1 vccd1 _15909_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_172_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17035_ _17035_/A _17035_/B vssd1 vssd1 vccd1 vccd1 _17035_/Y sky130_fd_sc_hd__nand2_1
XFILLER_7_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14247_ _14247_/A _14330_/B vssd1 vssd1 vccd1 vccd1 _14247_/Y sky130_fd_sc_hd__nor2_1
X_11459_ _11459_/A _11479_/B _12337_/S vssd1 vssd1 vccd1 vccd1 _11459_/X sky130_fd_sc_hd__and3_1
XFILLER_217_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14178_ _18695_/Q _13940_/X _13714_/X _18698_/Q vssd1 vssd1 vccd1 vccd1 _14178_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_217_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13129_ _13129_/A _18025_/Q vssd1 vssd1 vccd1 vccd1 _13130_/A sky130_fd_sc_hd__and2_1
XTAP_624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18986_ _18986_/CLK _18986_/D vssd1 vssd1 vccd1 vccd1 _18986_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17937_ _18204_/CLK _17937_/D vssd1 vssd1 vccd1 vccd1 _17937_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_152_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_213_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_1272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_213_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17868_ _19031_/CLK _17868_/D vssd1 vssd1 vccd1 vccd1 _17868_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_187_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19061__32 vssd1 vssd1 vccd1 vccd1 _19061__32/HI _19155_/A sky130_fd_sc_hd__conb_1
XFILLER_226_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16819_ _18136_/Q _17278_/B vssd1 vssd1 vccd1 vccd1 _16952_/A sky130_fd_sc_hd__nand2_1
XFILLER_38_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_187_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17799_ _17851_/CLK _17799_/D vssd1 vssd1 vccd1 vccd1 _17799_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_4_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_228_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_224_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09222_ _09222_/A _09222_/B vssd1 vssd1 vccd1 vccd1 _09222_/Y sky130_fd_sc_hd__nand2_1
XFILLER_22_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09153_ _09153_/A _09153_/B _10722_/A _09153_/D vssd1 vssd1 vccd1 vccd1 _09154_/C
+ sky130_fd_sc_hd__and4_1
XFILLER_72_1295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_120_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09084_ _09084_/A vssd1 vssd1 vccd1 vccd1 _19180_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_120_1238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09986_ _09986_/A vssd1 vssd1 vccd1 vccd1 _10955_/S sky130_fd_sc_hd__buf_4
XFILLER_104_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08937_ _08941_/A vssd1 vssd1 vccd1 vccd1 _08937_/Y sky130_fd_sc_hd__inv_2
XFILLER_44_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_218_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_218_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10830_ _09227_/C _09232_/B _09237_/D _09232_/D _10695_/A _10664_/A vssd1 vssd1 vccd1
+ vccd1 _10830_/X sky130_fd_sc_hd__mux4_2
XFILLER_164_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10761_ _10864_/A _10757_/B _10758_/X _10760_/X _10622_/Y vssd1 vssd1 vccd1 vccd1
+ _10761_/X sky130_fd_sc_hd__o311a_1
XFILLER_186_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_213_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12500_ _12498_/Y _12499_/X _12487_/Y vssd1 vssd1 vccd1 vccd1 _12500_/X sky130_fd_sc_hd__o21ba_1
XFILLER_9_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13480_ _13480_/A _13480_/B vssd1 vssd1 vccd1 vccd1 _18163_/D sky130_fd_sc_hd__nor2_1
X_10692_ _10757_/B vssd1 vssd1 vccd1 vccd1 _12094_/A sky130_fd_sc_hd__buf_2
XFILLER_164_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12431_ _12439_/A _12430_/B _12430_/C vssd1 vssd1 vccd1 vccd1 _12432_/C sky130_fd_sc_hd__a21o_1
XFILLER_12_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15150_ _15162_/A _15150_/B _15199_/C vssd1 vssd1 vccd1 vccd1 _15150_/X sky130_fd_sc_hd__or3_1
XFILLER_172_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12362_ _12387_/A vssd1 vssd1 vccd1 vccd1 _12467_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_181_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14101_ _18659_/Q _13617_/A _14099_/X _14100_/X vssd1 vssd1 vccd1 vccd1 _14101_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_148_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11313_ _11334_/A _11313_/B vssd1 vssd1 vccd1 vccd1 _11313_/X sky130_fd_sc_hd__and2b_1
X_15081_ _18395_/Q _18359_/Q _15081_/S vssd1 vssd1 vccd1 vccd1 _15081_/X sky130_fd_sc_hd__mux2_1
X_12293_ _12287_/Y _12293_/B _12313_/B vssd1 vssd1 vccd1 vccd1 _12294_/A sky130_fd_sc_hd__and3b_1
XFILLER_4_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14032_ _18251_/Q _13596_/X _13630_/X _18233_/Q vssd1 vssd1 vccd1 vccd1 _14032_/X
+ sky130_fd_sc_hd__a22o_1
X_11244_ _11244_/A vssd1 vssd1 vccd1 vccd1 _17823_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_175_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_180_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18840_ _18845_/CLK _18840_/D vssd1 vssd1 vccd1 vccd1 _18840_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_121_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11175_ _11175_/A vssd1 vssd1 vccd1 vccd1 _17805_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_68_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_132_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10126_ _10131_/A _10131_/B vssd1 vssd1 vccd1 vccd1 _10456_/A sky130_fd_sc_hd__xor2_4
X_18771_ _18799_/CLK _18771_/D vssd1 vssd1 vccd1 vccd1 _18771_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_122_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15983_ _18609_/Q _18573_/Q _15990_/S vssd1 vssd1 vccd1 vccd1 _15983_/X sky130_fd_sc_hd__mux2_1
XTAP_5651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17722_ _17722_/A vssd1 vssd1 vccd1 vccd1 _19005_/D sky130_fd_sc_hd__clkbuf_1
XTAP_5673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14934_ _18359_/Q _18323_/Q _14934_/S vssd1 vssd1 vccd1 vccd1 _14934_/X sky130_fd_sc_hd__mux2_1
X_10057_ _10055_/X _10056_/X _10956_/B vssd1 vssd1 vccd1 vccd1 _10057_/X sky130_fd_sc_hd__mux2_1
XTAP_5684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17653_ _17653_/A vssd1 vssd1 vccd1 vccd1 _18975_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_75_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_224_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14865_ _14977_/A vssd1 vssd1 vccd1 vccd1 _14958_/A sky130_fd_sc_hd__buf_2
XTAP_4994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_223_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16604_ _18756_/Q _18720_/Q _16617_/S vssd1 vssd1 vccd1 vccd1 _16604_/X sky130_fd_sc_hd__mux2_1
XFILLER_169_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13816_ _18939_/Q _13670_/X _13766_/A _18915_/Q vssd1 vssd1 vccd1 vccd1 _13816_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_17_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17584_ _17587_/A _17584_/B vssd1 vssd1 vccd1 vccd1 _17585_/A sky130_fd_sc_hd__and2_1
X_14796_ _14810_/A _14802_/B vssd1 vssd1 vccd1 vccd1 _14796_/Y sky130_fd_sc_hd__nand2_1
XFILLER_223_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16535_ _16572_/A _16538_/B vssd1 vssd1 vccd1 vccd1 _16535_/Y sky130_fd_sc_hd__nand2_1
X_13747_ _18336_/Q _13730_/X _13732_/X _18327_/Q _13746_/X vssd1 vssd1 vccd1 vccd1
+ _13747_/X sky130_fd_sc_hd__a221o_2
XFILLER_50_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10959_ _09711_/A _10954_/X _10958_/X _10010_/X vssd1 vssd1 vccd1 vccd1 _10959_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_44_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_188_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_189_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16466_ _16757_/A _16501_/B vssd1 vssd1 vccd1 vccd1 _16475_/B sky130_fd_sc_hd__nor2_2
XFILLER_176_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_231_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13678_ _18531_/Q _13489_/A _13763_/A _18546_/Q vssd1 vssd1 vccd1 vccd1 _13678_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_108_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18205_ _18991_/CLK _18205_/D vssd1 vssd1 vccd1 vccd1 _18205_/Q sky130_fd_sc_hd__dfxtp_1
X_15417_ _15445_/A _15417_/B vssd1 vssd1 vccd1 vccd1 _15417_/Y sky130_fd_sc_hd__nand2_1
XFILLER_31_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19185_ _19185_/A _09001_/Y vssd1 vssd1 vccd1 vccd1 io_out[23] sky130_fd_sc_hd__ebufn_8
X_12629_ _12629_/A vssd1 vssd1 vccd1 vccd1 _12630_/B sky130_fd_sc_hd__inv_2
X_16397_ _16434_/A _16692_/B _16422_/C vssd1 vssd1 vccd1 vccd1 _16397_/X sky130_fd_sc_hd__or3_1
XFILLER_157_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18136_ _18254_/CLK _18136_/D vssd1 vssd1 vccd1 vccd1 _18136_/Q sky130_fd_sc_hd__dfxtp_1
X_15348_ _18457_/Q _18421_/Q _15356_/S vssd1 vssd1 vccd1 vccd1 _15348_/X sky130_fd_sc_hd__mux2_1
XFILLER_89_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_117_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18067_ _18072_/CLK _18067_/D vssd1 vssd1 vccd1 vccd1 _18067_/Q sky130_fd_sc_hd__dfxtp_1
X_15279_ _15279_/A _15279_/B _15279_/C vssd1 vssd1 vccd1 vccd1 _15279_/X sky130_fd_sc_hd__or3_1
XFILLER_172_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17018_ _17032_/A _17023_/B vssd1 vssd1 vccd1 vccd1 _17018_/Y sky130_fd_sc_hd__nand2_1
XFILLER_104_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09840_ _09839_/A _09840_/B vssd1 vssd1 vccd1 vccd1 _09840_/X sky130_fd_sc_hd__and2b_1
XFILLER_113_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09771_ _09777_/A _09785_/B vssd1 vssd1 vccd1 vccd1 _09781_/B sky130_fd_sc_hd__xnor2_2
XFILLER_100_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18969_ _18972_/CLK _18969_/D vssd1 vssd1 vccd1 vccd1 _18969_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_227_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_226_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_215_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_226_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_2_2_0_wb_clk_i clkbuf_2_3_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_2_2_1_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_22_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_224_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_224_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09205_ _18692_/Q _18691_/Q _18690_/Q vssd1 vssd1 vccd1 vccd1 _09209_/A sky130_fd_sc_hd__or3_4
XFILLER_22_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09136_ _09136_/A _09136_/B _09136_/C _09136_/D vssd1 vssd1 vccd1 vccd1 _09137_/C
+ sky130_fd_sc_hd__and4_1
XFILLER_33_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_159_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09067_ _09072_/A _09069_/B _17827_/Q vssd1 vssd1 vccd1 vccd1 _09068_/A sky130_fd_sc_hd__and3_4
XFILLER_190_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_1306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09969_ _09969_/A vssd1 vssd1 vccd1 vccd1 _09969_/X sky130_fd_sc_hd__clkbuf_4
XTAP_4202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12980_ _12975_/A _12958_/B _12970_/A _12976_/B vssd1 vssd1 vccd1 vccd1 _12980_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_58_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11931_ _11951_/A _11951_/B _17792_/Q vssd1 vssd1 vccd1 vccd1 _11983_/B sky130_fd_sc_hd__o21ai_2
XTAP_3545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14650_ _16919_/A vssd1 vssd1 vccd1 vccd1 _15241_/A sky130_fd_sc_hd__buf_6
XFILLER_150_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11862_ _12257_/A vssd1 vssd1 vccd1 vccd1 _17764_/A sky130_fd_sc_hd__buf_4
XFILLER_72_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13601_ _18705_/Q _13577_/X _13590_/X _13600_/X vssd1 vssd1 vccd1 vccd1 _13601_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_150_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10813_ _10813_/A _10813_/B vssd1 vssd1 vccd1 vccd1 _10813_/X sky130_fd_sc_hd__or2_1
XTAP_2877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14581_ _14651_/A _15184_/A vssd1 vssd1 vccd1 vccd1 _14589_/B sky130_fd_sc_hd__nor2_1
XTAP_2888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11793_ _11740_/C _11789_/Y _11786_/Y _11749_/B _11792_/X vssd1 vssd1 vccd1 vccd1
+ _11793_/X sky130_fd_sc_hd__a221o_1
XTAP_2899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16320_ _18687_/Q _18651_/Q _16324_/S vssd1 vssd1 vccd1 vccd1 _16320_/X sky130_fd_sc_hd__mux2_1
XFILLER_159_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_186_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13532_ _13532_/A vssd1 vssd1 vccd1 vccd1 _13576_/A sky130_fd_sc_hd__buf_6
XFILLER_207_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10744_ _10664_/A _10741_/X _10743_/X _10805_/B vssd1 vssd1 vccd1 vccd1 _10744_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_213_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16251_ _16265_/A _16256_/B vssd1 vssd1 vccd1 vccd1 _16251_/Y sky130_fd_sc_hd__nand2_1
XFILLER_159_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13463_ _13467_/A _13463_/B vssd1 vssd1 vccd1 vccd1 _18155_/D sky130_fd_sc_hd__nor2_1
XFILLER_51_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10675_ _10675_/A _10820_/B vssd1 vssd1 vccd1 vccd1 _12101_/A sky130_fd_sc_hd__xnor2_4
X_15202_ _18424_/Q _18388_/Q _15226_/S vssd1 vssd1 vccd1 vccd1 _15202_/X sky130_fd_sc_hd__mux2_1
XFILLER_167_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12414_ _12414_/A _12414_/B _12414_/C vssd1 vssd1 vccd1 vccd1 _12415_/B sky130_fd_sc_hd__or3_1
X_16182_ _16188_/B _16179_/X _16181_/X _16162_/X vssd1 vssd1 vccd1 vccd1 _18618_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_16_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13394_ _13375_/A _17996_/Q _17997_/Q _13394_/D vssd1 vssd1 vccd1 vccd1 _13405_/B
+ sky130_fd_sc_hd__and4bb_4
XFILLER_12_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15133_ _15132_/B _15130_/X _15132_/Y _15123_/X vssd1 vssd1 vccd1 vccd1 _18371_/D
+ sky130_fd_sc_hd__o211a_1
X_12345_ _11463_/B _12336_/X _12328_/B _17888_/Q vssd1 vssd1 vccd1 vccd1 _12346_/C
+ sky130_fd_sc_hd__o211a_1
XFILLER_103_1277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15064_ _15064_/A vssd1 vssd1 vccd1 vccd1 _15112_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_138_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12276_ _17869_/Q _13066_/B _12276_/C vssd1 vssd1 vccd1 vccd1 _12277_/A sky130_fd_sc_hd__and3_1
XFILLER_107_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_218_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14015_ _14015_/A vssd1 vssd1 vccd1 vccd1 _14015_/X sky130_fd_sc_hd__buf_4
X_11227_ _11232_/C _11227_/B _11243_/A vssd1 vssd1 vccd1 vccd1 _11228_/A sky130_fd_sc_hd__and3b_1
XFILLER_229_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_214_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18823_ _18823_/CLK _18823_/D vssd1 vssd1 vccd1 vccd1 _18823_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_95_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11158_ _11501_/A vssd1 vssd1 vccd1 vccd1 _11780_/A sky130_fd_sc_hd__clkbuf_2
Xclkbuf_leaf_156_wb_clk_i _18102_/CLK vssd1 vssd1 vccd1 vccd1 _19028_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_96_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10109_ _10069_/X _10081_/X _10108_/X _10966_/B vssd1 vssd1 vccd1 vccd1 _10109_/X
+ sky130_fd_sc_hd__a22o_1
X_15966_ _16014_/A vssd1 vssd1 vccd1 vccd1 _15990_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_191_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18754_ _18788_/CLK _18754_/D vssd1 vssd1 vccd1 vccd1 _18754_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_49_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11089_ _17792_/Q vssd1 vssd1 vccd1 vccd1 _11963_/A sky130_fd_sc_hd__clkbuf_2
XTAP_5470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14917_ _15527_/A _14989_/C vssd1 vssd1 vccd1 vccd1 _14924_/B sky130_fd_sc_hd__nor2_2
X_17705_ _12373_/A _17704_/Y _17705_/S vssd1 vssd1 vccd1 vccd1 _17706_/A sky130_fd_sc_hd__mux2_1
XFILLER_36_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18685_ _18686_/CLK _18685_/D vssd1 vssd1 vccd1 vccd1 _18685_/Q sky130_fd_sc_hd__dfxtp_2
X_15897_ _15938_/A _15900_/B vssd1 vssd1 vccd1 vccd1 _15897_/Y sky130_fd_sc_hd__nand2_1
XTAP_4780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_223_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14848_ _18338_/Q _18302_/Q _14848_/S vssd1 vssd1 vccd1 vccd1 _14848_/X sky130_fd_sc_hd__mux2_1
X_17636_ _17635_/Y _17604_/X _17591_/X vssd1 vssd1 vccd1 vccd1 _17636_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_36_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17567_ _18183_/Q vssd1 vssd1 vccd1 vccd1 _17567_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_225_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14779_ _18284_/Q _14777_/B _14777_/Y _14778_/X vssd1 vssd1 vccd1 vccd1 _18284_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_90_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16518_ _16555_/A _16666_/B _16568_/C vssd1 vssd1 vccd1 vccd1 _16518_/X sky130_fd_sc_hd__or3_1
XFILLER_225_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17498_ _17501_/B _17495_/X _17496_/Y _17497_/X vssd1 vssd1 vccd1 vccd1 _18937_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_220_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16449_ _18719_/Q _18683_/Q _16449_/S vssd1 vssd1 vccd1 vccd1 _16449_/X sky130_fd_sc_hd__mux2_1
XFILLER_143_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19237_ _19237_/A _08940_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[37] sky130_fd_sc_hd__ebufn_8
XFILLER_34_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19168_ _19168_/A _09015_/Y vssd1 vssd1 vccd1 vccd1 io_out[6] sky130_fd_sc_hd__ebufn_8
XFILLER_219_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_1366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18119_ _18125_/CLK _18119_/D vssd1 vssd1 vccd1 vccd1 _18119_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_145_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09823_ _18126_/Q _09844_/A vssd1 vssd1 vccd1 vccd1 _12112_/A sky130_fd_sc_hd__or2_1
XFILLER_101_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09754_ _17783_/Q vssd1 vssd1 vccd1 vccd1 _09784_/A sky130_fd_sc_hd__inv_2
XFILLER_41_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_227_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_227_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09685_ _09704_/A _09704_/B vssd1 vssd1 vccd1 vccd1 _09991_/A sky130_fd_sc_hd__nor2_2
XFILLER_54_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_1290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_223_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_210_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_168_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_196_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_202_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_211_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10460_ _10547_/B _10419_/A _10455_/X _10459_/X vssd1 vssd1 vccd1 vccd1 _10460_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_148_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09119_ _09119_/A _09119_/B _09119_/C _10350_/A vssd1 vssd1 vccd1 vccd1 _09120_/C
+ sky130_fd_sc_hd__and4_1
X_10391_ _10391_/A _10391_/B vssd1 vssd1 vccd1 vccd1 _10391_/X sky130_fd_sc_hd__or2_1
XFILLER_11_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12130_ _12130_/A _13649_/B vssd1 vssd1 vccd1 vccd1 _12132_/C sky130_fd_sc_hd__xnor2_1
XFILLER_89_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12061_ _12061_/A _12126_/B vssd1 vssd1 vccd1 vccd1 _12061_/X sky130_fd_sc_hd__xor2_1
XFILLER_78_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11012_ _11012_/A vssd1 vssd1 vccd1 vccd1 _19174_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_150_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15820_ _16287_/A _15894_/C vssd1 vssd1 vccd1 vccd1 _15829_/B sky130_fd_sc_hd__nor2_1
XTAP_4010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_219_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_218_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15751_ _15751_/A _15754_/B vssd1 vssd1 vccd1 vccd1 _15751_/Y sky130_fd_sc_hd__nand2_1
XTAP_3320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_60 _11896_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12963_ _17984_/Q _12955_/X _12960_/X _12962_/Y _12949_/Y vssd1 vssd1 vccd1 vccd1
+ _12963_/X sky130_fd_sc_hd__a221o_1
XFILLER_79_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_71 _13529_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14702_ _14702_/A vssd1 vssd1 vccd1 vccd1 _16219_/A sky130_fd_sc_hd__buf_6
XTAP_4098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_82 _13591_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_218_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_205_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18470_ _18473_/CLK _18470_/D vssd1 vssd1 vccd1 vccd1 _18470_/Q sky130_fd_sc_hd__dfxtp_2
XINSDIODE2_93 _13677_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11914_ _18128_/Q _10256_/A _11913_/X vssd1 vssd1 vccd1 vccd1 _11915_/B sky130_fd_sc_hd__a21bo_1
X_15682_ _18499_/Q _15683_/B _15680_/Y _15681_/X vssd1 vssd1 vccd1 vccd1 _18499_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_2630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12894_ _12792_/X _12895_/C _12893_/Y vssd1 vssd1 vccd1 vccd1 _17961_/D sky130_fd_sc_hd__a21oi_1
XTAP_3386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17421_ _17497_/A vssd1 vssd1 vccd1 vccd1 _17421_/X sky130_fd_sc_hd__buf_2
XTAP_2652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14633_ _18250_/Q _14635_/B _14632_/Y _14629_/X vssd1 vssd1 vccd1 vccd1 _18250_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_72_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11845_ _11845_/A _11845_/B _11845_/C vssd1 vssd1 vccd1 vccd1 _11850_/B sky130_fd_sc_hd__and3_1
XFILLER_45_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_202_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17352_ _17370_/A vssd1 vssd1 vccd1 vccd1 _17367_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_207_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_198_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14564_ _14672_/A vssd1 vssd1 vccd1 vccd1 _17674_/A sky130_fd_sc_hd__buf_2
X_11776_ _11780_/A _11776_/B vssd1 vssd1 vccd1 vccd1 _11776_/Y sky130_fd_sc_hd__xnor2_1
XTAP_1984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16303_ _16305_/B _16301_/X _16302_/Y _16295_/X vssd1 vssd1 vccd1 vccd1 _18646_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_207_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13515_ _13515_/A vssd1 vssd1 vccd1 vccd1 _13515_/X sky130_fd_sc_hd__buf_6
XFILLER_18_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10727_ _09114_/A _09119_/B _10841_/A vssd1 vssd1 vccd1 vccd1 _10727_/X sky130_fd_sc_hd__mux2_1
X_17283_ _17304_/A vssd1 vssd1 vccd1 vccd1 _17283_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_202_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14495_ _14495_/A vssd1 vssd1 vccd1 vccd1 _18221_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_201_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19022_ _19026_/CLK _19022_/D vssd1 vssd1 vccd1 vccd1 _19022_/Q sky130_fd_sc_hd__dfxtp_1
X_16234_ _16348_/A vssd1 vssd1 vccd1 vccd1 _16327_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_186_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13446_ _13446_/A _13452_/A vssd1 vssd1 vccd1 vccd1 _13446_/Y sky130_fd_sc_hd__nor2_1
X_10658_ _10813_/B vssd1 vssd1 vccd1 vccd1 _10812_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_16_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16165_ _16757_/A _16205_/B vssd1 vssd1 vccd1 vccd1 _16175_/B sky130_fd_sc_hd__nor2_2
XFILLER_115_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13377_ _09752_/A _13344_/X _13337_/X _13379_/B vssd1 vssd1 vccd1 vccd1 _18111_/D
+ sky130_fd_sc_hd__o211a_1
X_10589_ _09332_/B _09327_/B _09337_/C _09327_/C _10089_/S _10036_/X vssd1 vssd1 vccd1
+ vccd1 _10589_/X sky130_fd_sc_hd__mux4_2
XFILLER_6_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15116_ _15118_/B _15114_/X _15115_/Y _15103_/X vssd1 vssd1 vccd1 vccd1 _18367_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_142_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12328_ _13418_/C _12328_/B vssd1 vssd1 vccd1 vccd1 _12347_/B sky130_fd_sc_hd__nor2_2
X_16096_ _16132_/A _16096_/B vssd1 vssd1 vccd1 vccd1 _16096_/Y sky130_fd_sc_hd__nand2_1
XFILLER_181_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15047_ _15049_/B _15044_/X _15045_/Y _15046_/X vssd1 vssd1 vccd1 vccd1 _18349_/D
+ sky130_fd_sc_hd__o211a_1
X_12259_ _12259_/A vssd1 vssd1 vccd1 vccd1 _17864_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_69_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_218_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_1367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_205_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18806_ _18806_/CLK _18806_/D vssd1 vssd1 vccd1 vccd1 _18806_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_83_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16998_ _17035_/A _16998_/B vssd1 vssd1 vccd1 vccd1 _16998_/Y sky130_fd_sc_hd__nand2_1
XFILLER_55_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18737_ _18765_/CLK _18737_/D vssd1 vssd1 vccd1 vccd1 _18737_/Q sky130_fd_sc_hd__dfxtp_1
X_15949_ _15960_/B _15945_/X _15946_/X _15948_/X vssd1 vssd1 vccd1 vccd1 _18564_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_83_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_225_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09470_ _09470_/A _09474_/A vssd1 vssd1 vccd1 vccd1 _09471_/B sky130_fd_sc_hd__and2_1
XFILLER_224_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18668_ _18668_/CLK _18668_/D vssd1 vssd1 vccd1 vccd1 _18668_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_149_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_221_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17619_ _17616_/Y _17552_/X _18967_/Q vssd1 vssd1 vccd1 vccd1 _17619_/X sky130_fd_sc_hd__a21o_1
XFILLER_224_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18599_ _18608_/CLK _18599_/D vssd1 vssd1 vccd1 vccd1 _18599_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_211_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_225_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_53_wb_clk_i clkbuf_5_16_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18785_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_211_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_1327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_220_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_1264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_191_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_69_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_219_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09806_ _09806_/A _09806_/B vssd1 vssd1 vccd1 vccd1 _09807_/B sky130_fd_sc_hd__xnor2_1
XFILLER_75_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_219_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_216_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09737_ _09739_/B _09739_/A vssd1 vssd1 vccd1 vccd1 _09748_/A sky130_fd_sc_hd__or2b_1
XFILLER_41_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_1292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09668_ _09668_/A _09668_/B vssd1 vssd1 vccd1 vccd1 _12070_/A sky130_fd_sc_hd__xnor2_4
XFILLER_83_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_227_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_1366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_203_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_188_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_231_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09599_ _09600_/A _09600_/B _09600_/C vssd1 vssd1 vccd1 vccd1 _09601_/A sky130_fd_sc_hd__nor3_1
XFILLER_199_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11630_ _12221_/A _11617_/X _11628_/Y _11609_/X _11629_/Y vssd1 vssd1 vccd1 vccd1
+ _11630_/X sky130_fd_sc_hd__o32a_1
XTAP_1269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_230_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11561_ _17868_/Q vssd1 vssd1 vccd1 vccd1 _11563_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_10_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13300_ _18042_/Q _18045_/Q _18044_/Q _18047_/Q vssd1 vssd1 vccd1 vccd1 _13303_/A
+ sky130_fd_sc_hd__or4_1
XFILLER_155_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10512_ _10926_/A _10512_/B _10512_/C vssd1 vssd1 vccd1 vccd1 _10512_/X sky130_fd_sc_hd__and3_1
XFILLER_195_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14280_ _14224_/Y _14335_/B _14355_/B vssd1 vssd1 vccd1 vccd1 _14280_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_156_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11492_ _17890_/Q _11485_/X _11488_/Y _11490_/Y _11491_/Y vssd1 vssd1 vccd1 vccd1
+ _11492_/X sky130_fd_sc_hd__a41o_1
XFILLER_10_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13231_ _13233_/A _18071_/Q vssd1 vssd1 vccd1 vccd1 _13232_/A sky130_fd_sc_hd__and2_1
XFILLER_10_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10443_ _10443_/A vssd1 vssd1 vccd1 vccd1 _10443_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_171_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_1323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_1334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13162_ _13164_/A _18040_/Q vssd1 vssd1 vccd1 vccd1 _13163_/A sky130_fd_sc_hd__and2_1
XFILLER_40_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10374_ _10598_/A _10374_/B vssd1 vssd1 vccd1 vccd1 _10374_/X sky130_fd_sc_hd__or2_1
XFILLER_174_1326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12113_ _09843_/A _12112_/A _09833_/B _12111_/Y _12112_/X vssd1 vssd1 vccd1 vccd1
+ _12117_/A sky130_fd_sc_hd__a311o_1
XFILLER_215_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_1359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13093_ _13093_/A vssd1 vssd1 vccd1 vccd1 _18008_/D sky130_fd_sc_hd__clkbuf_1
X_17970_ _18108_/CLK _17970_/D vssd1 vssd1 vccd1 vccd1 _17970_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_46_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16921_ _18831_/Q _18795_/Q _16925_/S vssd1 vssd1 vccd1 vccd1 _16921_/X sky130_fd_sc_hd__mux2_1
X_12044_ _12044_/A _13693_/A vssd1 vssd1 vccd1 vccd1 _12101_/B sky130_fd_sc_hd__nand2_2
XFILLER_215_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16852_ _18816_/Q _18780_/Q _16864_/S vssd1 vssd1 vccd1 vccd1 _16852_/X sky130_fd_sc_hd__mux2_1
XFILLER_65_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_226_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_120_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15803_ _15823_/A vssd1 vssd1 vccd1 vccd1 _15803_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_133_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16783_ _16783_/A _16794_/B vssd1 vssd1 vccd1 vccd1 _16792_/B sky130_fd_sc_hd__nor2_1
X_13995_ _18559_/Q _13677_/X _13721_/A _18583_/Q vssd1 vssd1 vccd1 vccd1 _13995_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_18_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18522_ _18532_/CLK _18522_/D vssd1 vssd1 vccd1 vccd1 _18522_/Q sky130_fd_sc_hd__dfxtp_2
X_15734_ _15734_/A _16032_/B _15748_/C vssd1 vssd1 vccd1 vccd1 _15734_/X sky130_fd_sc_hd__or3_1
XFILLER_19_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12946_ _12946_/A vssd1 vssd1 vccd1 vccd1 _12961_/A sky130_fd_sc_hd__clkbuf_2
XTAP_3150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18453_ _18458_/CLK _18453_/D vssd1 vssd1 vccd1 vccd1 _18453_/Q sky130_fd_sc_hd__dfxtp_2
X_15665_ _18531_/Q _18495_/Q _15665_/S vssd1 vssd1 vccd1 vccd1 _15665_/X sky130_fd_sc_hd__mux2_1
XFILLER_209_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_206_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_181_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12877_ _17955_/Q _17956_/Q _12877_/C vssd1 vssd1 vccd1 vccd1 _12881_/B sky130_fd_sc_hd__and3_1
XTAP_2460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14616_ _14357_/X _14608_/X _14612_/X _14615_/Y _11822_/X vssd1 vssd1 vccd1 vccd1
+ _18247_/D sky130_fd_sc_hd__o311a_1
XFILLER_33_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17404_ _17453_/A _17408_/B vssd1 vssd1 vccd1 vccd1 _17404_/Y sky130_fd_sc_hd__nand2_1
X_18384_ _18387_/CLK _18384_/D vssd1 vssd1 vccd1 vccd1 _18384_/Q sky130_fd_sc_hd__dfxtp_4
X_11828_ _11828_/A _11828_/B vssd1 vssd1 vccd1 vccd1 _11828_/Y sky130_fd_sc_hd__nand2_2
X_15596_ _15594_/B _15593_/X _15594_/Y _15595_/X vssd1 vssd1 vccd1 vccd1 _18479_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_1770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17335_ _18895_/Q _17336_/B _17334_/Y _17324_/X vssd1 vssd1 vccd1 vccd1 _18895_/D
+ sky130_fd_sc_hd__o211a_1
X_14547_ _14593_/A vssd1 vssd1 vccd1 vccd1 _17602_/A sky130_fd_sc_hd__buf_2
XFILLER_230_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11759_ _11767_/C vssd1 vssd1 vccd1 vccd1 _11761_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_197_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17266_ _17331_/A vssd1 vssd1 vccd1 vccd1 _17399_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_201_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14478_ _18214_/Q _14480_/B vssd1 vssd1 vccd1 vccd1 _14479_/A sky130_fd_sc_hd__and2_1
XFILLER_174_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16217_ _16268_/A _16217_/B vssd1 vssd1 vccd1 vccd1 _16217_/Y sky130_fd_sc_hd__nand2_1
X_19005_ _19009_/CLK _19005_/D vssd1 vssd1 vccd1 vccd1 _19005_/Q sky130_fd_sc_hd__dfxtp_1
X_13429_ _13429_/A vssd1 vssd1 vccd1 vccd1 _13429_/Y sky130_fd_sc_hd__inv_2
XFILLER_60_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17197_ _17197_/A vssd1 vssd1 vccd1 vccd1 _17197_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_16148_ _16147_/B _16145_/X _16147_/Y _16139_/X vssd1 vssd1 vccd1 vccd1 _18611_/D
+ sky130_fd_sc_hd__o211a_1
Xclkbuf_leaf_171_wb_clk_i clkbuf_5_11_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18044_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_143_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16079_ _16082_/B _16076_/X _16078_/Y _16074_/X vssd1 vssd1 vccd1 vccd1 _18595_/D
+ sky130_fd_sc_hd__o211a_1
Xclkbuf_leaf_100_wb_clk_i clkbuf_5_28_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18511_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_130_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08970_ _08972_/A vssd1 vssd1 vccd1 vccd1 _08970_/Y sky130_fd_sc_hd__inv_2
XFILLER_9_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_216_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_229_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_229_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput1 active vssd1 vssd1 vccd1 vccd1 input1/X sky130_fd_sc_hd__buf_12
XFILLER_151_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09522_ _14332_/S vssd1 vssd1 vccd1 vccd1 _14267_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_25_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_225_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09453_ _09430_/C _09430_/D _09452_/X _09138_/A vssd1 vssd1 vccd1 vccd1 _09454_/C
+ sky130_fd_sc_hd__a31o_1
XFILLER_80_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_212_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09384_ _18377_/Q _18376_/Q _18375_/Q vssd1 vssd1 vccd1 vccd1 _09972_/A sky130_fd_sc_hd__or3_4
XFILLER_101_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_221_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_177_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_193_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10090_ _10088_/X _10089_/X _10090_/S vssd1 vssd1 vccd1 vccd1 _10090_/X sky130_fd_sc_hd__mux2_1
XFILLER_86_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12800_ _12597_/B _17953_/Q _12871_/A _12609_/B vssd1 vssd1 vccd1 vccd1 _12800_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_90_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13780_ _13780_/A vssd1 vssd1 vccd1 vccd1 _13780_/X sky130_fd_sc_hd__buf_8
XFILLER_27_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10992_ _10985_/X _09523_/X _10977_/X _10982_/A _14204_/B vssd1 vssd1 vccd1 vccd1
+ _18996_/D sky130_fd_sc_hd__a32o_1
XFILLER_210_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_231_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12731_ _12919_/B vssd1 vssd1 vccd1 vccd1 _13310_/A sky130_fd_sc_hd__buf_2
XFILLER_16_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_163_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_231_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15450_ _16962_/A vssd1 vssd1 vccd1 vccd1 _16043_/B sky130_fd_sc_hd__buf_2
XFILLER_31_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_203_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12662_ _12662_/A _12662_/B vssd1 vssd1 vccd1 vccd1 _12663_/B sky130_fd_sc_hd__nor2_1
XFILLER_230_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_231_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14401_ _14428_/A vssd1 vssd1 vccd1 vccd1 _14401_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_204_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_180_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11613_ _11624_/B vssd1 vssd1 vccd1 vccd1 _12221_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_230_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15381_ _15423_/A _15984_/B _15423_/C vssd1 vssd1 vccd1 vccd1 _15381_/X sky130_fd_sc_hd__or3_1
XFILLER_204_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_212_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12593_ _17923_/Q _12569_/X _12590_/Y _12592_/X _12548_/X vssd1 vssd1 vccd1 vccd1
+ _17923_/D sky130_fd_sc_hd__a221o_1
XFILLER_204_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17120_ _17120_/A _17549_/B vssd1 vssd1 vccd1 vccd1 _17184_/A sky130_fd_sc_hd__or2_2
X_14332_ _14331_/X _10605_/A _14332_/S vssd1 vssd1 vccd1 vccd1 _14334_/B sky130_fd_sc_hd__mux2_1
XFILLER_168_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11544_ _13526_/A vssd1 vssd1 vccd1 vccd1 _12089_/B sky130_fd_sc_hd__buf_6
XFILLER_7_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_195_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17051_ _17056_/B _17049_/X _17050_/X _17040_/X vssd1 vssd1 vccd1 vccd1 _18825_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_7_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14263_ _14243_/X _14227_/X _14229_/X _14244_/X _18172_/Q vssd1 vssd1 vccd1 vccd1
+ _14263_/X sky130_fd_sc_hd__a311o_1
XFILLER_171_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11475_ _11478_/A _11472_/A _11463_/B _11377_/A vssd1 vssd1 vccd1 vccd1 _11475_/X
+ sky130_fd_sc_hd__a211o_1
X_16002_ _18614_/Q _18578_/Q _16010_/S vssd1 vssd1 vccd1 vccd1 _16002_/X sky130_fd_sc_hd__mux2_1
X_13214_ _13222_/A _18063_/Q vssd1 vssd1 vccd1 vccd1 _13215_/A sky130_fd_sc_hd__and2_1
X_10426_ _09136_/B _09126_/D _09126_/A _09131_/A _10235_/A _10413_/A vssd1 vssd1 vccd1
+ vccd1 _10427_/B sky130_fd_sc_hd__mux4_2
XFILLER_124_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14194_ _18226_/Q _18225_/Q _18224_/Q _18223_/Q vssd1 vssd1 vccd1 vccd1 _14196_/B
+ sky130_fd_sc_hd__or4_1
XFILLER_152_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13145_ _13151_/A _18032_/Q vssd1 vssd1 vccd1 vccd1 _13146_/A sky130_fd_sc_hd__and2_1
XFILLER_48_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10357_ _14260_/B _10354_/X _10356_/X _10338_/A vssd1 vssd1 vccd1 vccd1 _10357_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_140_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13076_ _18007_/Q _18009_/Q vssd1 vssd1 vccd1 vccd1 _13076_/X sky130_fd_sc_hd__xor2_1
X_17953_ _17959_/CLK _17953_/D vssd1 vssd1 vccd1 vccd1 _17953_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_140_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10288_ _10288_/A _10288_/B vssd1 vssd1 vccd1 vccd1 _10288_/Y sky130_fd_sc_hd__nor2_1
XFILLER_105_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16904_ _16903_/B _16900_/X _16903_/Y _16893_/X vssd1 vssd1 vccd1 vccd1 _18791_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_61_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12027_ _12027_/A _12027_/B _12027_/C _12027_/D vssd1 vssd1 vccd1 vccd1 _12028_/C
+ sky130_fd_sc_hd__or4_1
XFILLER_215_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17884_ _17884_/CLK _17884_/D vssd1 vssd1 vccd1 vccd1 _17884_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16835_ _16835_/A vssd1 vssd1 vccd1 vccd1 _17435_/A sky130_fd_sc_hd__buf_4
XFILLER_226_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_226_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13978_ _18352_/Q _13489_/A _13763_/A _18367_/Q vssd1 vssd1 vccd1 vccd1 _13978_/X
+ sky130_fd_sc_hd__a22o_1
X_16766_ _16766_/A vssd1 vssd1 vccd1 vccd1 _16784_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_207_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18505_ _18506_/CLK _18505_/D vssd1 vssd1 vccd1 vccd1 _18505_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_20_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15717_ _15717_/A vssd1 vssd1 vccd1 vccd1 _15733_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_146_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12929_ _12947_/A _12923_/Y _12928_/X _12760_/X vssd1 vssd1 vccd1 vccd1 _12930_/A
+ sky130_fd_sc_hd__o211a_1
X_16697_ _16766_/A vssd1 vssd1 vccd1 vccd1 _16715_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_185_1274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_222_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18436_ _18443_/CLK _18436_/D vssd1 vssd1 vccd1 vccd1 _18436_/Q sky130_fd_sc_hd__dfxtp_2
X_15648_ _18527_/Q _18491_/Q _15665_/S vssd1 vssd1 vccd1 vccd1 _15648_/X sky130_fd_sc_hd__mux2_1
XTAP_2290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15579_ _15630_/A _15583_/B vssd1 vssd1 vccd1 vccd1 _15579_/Y sky130_fd_sc_hd__nand2_1
X_18367_ _18367_/CLK _18367_/D vssd1 vssd1 vccd1 vccd1 _18367_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_187_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_222_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_187_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17318_ _17318_/A _17460_/B _17318_/C vssd1 vssd1 vccd1 vccd1 _17318_/X sky130_fd_sc_hd__or3_1
XFILLER_179_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18298_ _18308_/CLK _18298_/D vssd1 vssd1 vccd1 vccd1 _18298_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17249_ _17273_/A _17252_/B vssd1 vssd1 vccd1 vccd1 _17249_/Y sky130_fd_sc_hd__nand2_1
XFILLER_174_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_190_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_227_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_1310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08953_ _08954_/A vssd1 vssd1 vccd1 vccd1 _08953_/Y sky130_fd_sc_hd__inv_2
XTAP_4609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_229_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_186_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09505_ _18204_/Q _09505_/B vssd1 vssd1 vccd1 vccd1 _09506_/B sky130_fd_sc_hd__or2_1
XFILLER_225_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_213_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_1306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_1366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09436_ _09421_/A _09222_/Y _09454_/B _09432_/B vssd1 vssd1 vccd1 vccd1 _09474_/A
+ sky130_fd_sc_hd__o211a_2
XPHY_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_227_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_212_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09367_ _18269_/Q _18268_/Q _18267_/Q vssd1 vssd1 vccd1 vccd1 _09370_/B sky130_fd_sc_hd__or3_2
XFILLER_166_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09298_ _18509_/Q _18508_/Q _18507_/Q vssd1 vssd1 vccd1 vccd1 _09299_/D sky130_fd_sc_hd__or3_4
XFILLER_166_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11260_ _17799_/Q _17798_/Q vssd1 vssd1 vccd1 vccd1 _11287_/A sky130_fd_sc_hd__or2_1
XFILLER_106_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10211_ _10211_/A _10211_/B vssd1 vssd1 vccd1 vccd1 _10238_/A sky130_fd_sc_hd__nor2_2
X_11191_ _11210_/A _11191_/B _11193_/B vssd1 vssd1 vccd1 vccd1 _11192_/A sky130_fd_sc_hd__and3_1
XFILLER_122_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10142_ _10142_/A _10142_/B vssd1 vssd1 vccd1 vccd1 _10142_/Y sky130_fd_sc_hd__nor2_1
XFILLER_97_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14950_ _14949_/B _14947_/X _14949_/Y _14941_/X vssd1 vssd1 vccd1 vccd1 _18326_/D
+ sky130_fd_sc_hd__o211a_1
X_10073_ _10071_/X _10072_/X _10076_/S vssd1 vssd1 vccd1 vccd1 _10073_/X sky130_fd_sc_hd__mux2_1
XFILLER_212_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13901_ _18550_/Q _13663_/X _13664_/X _18526_/Q _13900_/X vssd1 vssd1 vccd1 vccd1
+ _13901_/X sky130_fd_sc_hd__a221o_1
XTAP_5888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14881_ _14881_/A vssd1 vssd1 vccd1 vccd1 _14881_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_87_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16620_ _16623_/B _16617_/X _16618_/Y _16619_/X vssd1 vssd1 vccd1 vccd1 _18724_/D
+ sky130_fd_sc_hd__o211a_1
X_13832_ _17709_/A _13832_/B vssd1 vssd1 vccd1 vccd1 _13833_/A sky130_fd_sc_hd__or2_1
XFILLER_21_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_223_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_204_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16551_ _16575_/A _16551_/B vssd1 vssd1 vccd1 vccd1 _16551_/Y sky130_fd_sc_hd__nand2_1
XINSDIODE2_207 _13492_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_218 _13785_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13763_ _13763_/A vssd1 vssd1 vccd1 vccd1 _13764_/A sky130_fd_sc_hd__buf_6
XFILLER_16_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XINSDIODE2_229 _15229_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10975_ _14282_/A vssd1 vssd1 vccd1 vccd1 _14272_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_90_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15502_ _15944_/A _15548_/B vssd1 vssd1 vccd1 vccd1 _15511_/B sky130_fd_sc_hd__nor2_2
X_12714_ _17940_/Q _18000_/Q vssd1 vssd1 vccd1 vccd1 _12748_/A sky130_fd_sc_hd__or2b_1
X_16482_ _16487_/B _16480_/X _16481_/X _16477_/X vssd1 vssd1 vccd1 vccd1 _18690_/D
+ sky130_fd_sc_hd__o211a_1
X_13694_ _13686_/X _13692_/X _13693_/Y vssd1 vssd1 vccd1 vccd1 _13694_/X sky130_fd_sc_hd__o21a_1
XFILLER_15_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15433_ _16949_/A vssd1 vssd1 vccd1 vccd1 _16030_/A sky130_fd_sc_hd__clkbuf_4
X_18221_ _18222_/CLK _18221_/D vssd1 vssd1 vccd1 vccd1 _18221_/Q sky130_fd_sc_hd__dfxtp_1
X_12645_ _12646_/A _12646_/B vssd1 vssd1 vccd1 vccd1 _12647_/A sky130_fd_sc_hd__and2_1
XFILLER_169_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_1280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15364_ _15366_/B _15361_/X _15362_/Y _15363_/X vssd1 vssd1 vccd1 vccd1 _18424_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_168_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18152_ _18997_/CLK _18152_/D vssd1 vssd1 vccd1 vccd1 _18152_/Q sky130_fd_sc_hd__dfxtp_2
X_12576_ _12561_/Y _12571_/X _12575_/Y vssd1 vssd1 vccd1 vccd1 _12576_/X sky130_fd_sc_hd__a21o_1
XFILLER_180_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_1204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17103_ _18875_/Q _18839_/Q _17114_/S vssd1 vssd1 vccd1 vccd1 _17103_/X sky130_fd_sc_hd__mux2_1
XFILLER_50_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14315_ _14299_/X _14282_/X _14283_/X _14300_/X _15903_/C vssd1 vssd1 vccd1 vccd1
+ _14315_/X sky130_fd_sc_hd__a311o_1
XFILLER_102_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11527_ _17873_/Q _11524_/X _11526_/X vssd1 vssd1 vccd1 vccd1 _11527_/Y sky130_fd_sc_hd__o21ai_1
X_18083_ _18087_/CLK _18083_/D vssd1 vssd1 vccd1 vccd1 _18083_/Q sky130_fd_sc_hd__dfxtp_1
X_15295_ _15562_/A vssd1 vssd1 vccd1 vccd1 _15358_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_156_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17034_ _18857_/Q _18821_/Q _17055_/S vssd1 vssd1 vccd1 vccd1 _17034_/X sky130_fd_sc_hd__mux2_1
XFILLER_176_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14246_ _14202_/X _14242_/X _14245_/X _13334_/X vssd1 vssd1 vccd1 vccd1 _18170_/D
+ sky130_fd_sc_hd__o211a_1
X_11458_ _17885_/Q vssd1 vssd1 vccd1 vccd1 _12337_/S sky130_fd_sc_hd__inv_2
XFILLER_109_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10409_ _10936_/S vssd1 vssd1 vccd1 vccd1 _12039_/A sky130_fd_sc_hd__clkbuf_4
X_14177_ _18686_/Q _13562_/A _13568_/A _18680_/Q _14176_/X vssd1 vssd1 vccd1 vccd1
+ _14177_/X sky130_fd_sc_hd__a221o_1
Xclkbuf_3_4_0_wb_clk_i clkbuf_3_5_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_4_9_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_125_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11389_ _11828_/A vssd1 vssd1 vccd1 vccd1 _11390_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_139_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13128_ _13128_/A vssd1 vssd1 vccd1 vccd1 _18023_/D sky130_fd_sc_hd__clkbuf_1
XTAP_614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18985_ _18986_/CLK _18985_/D vssd1 vssd1 vccd1 vccd1 _18985_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13059_ _13080_/A _13055_/B _13058_/B vssd1 vssd1 vccd1 vccd1 _13059_/Y sky130_fd_sc_hd__a21oi_1
X_17936_ _18204_/CLK _17936_/D vssd1 vssd1 vccd1 vccd1 _17936_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_100_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17867_ _19031_/CLK _17867_/D vssd1 vssd1 vccd1 vccd1 _17867_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_93_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_213_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_187_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16818_ _17423_/A _16963_/C vssd1 vssd1 vccd1 vccd1 _16833_/B sky130_fd_sc_hd__nor2_2
XFILLER_19_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17798_ _17851_/CLK _17798_/D vssd1 vssd1 vccd1 vccd1 _17798_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_187_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16749_ _16796_/A _16749_/B _16773_/C vssd1 vssd1 vccd1 vccd1 _16749_/X sky130_fd_sc_hd__or3_1
XFILLER_35_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_222_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_222_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09221_ _09188_/X _09221_/B _09430_/D vssd1 vssd1 vccd1 vccd1 _09222_/B sky130_fd_sc_hd__and3b_1
XFILLER_21_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18419_ _18423_/CLK _18419_/D vssd1 vssd1 vccd1 vccd1 _18419_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_61_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_222_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_148_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09152_ _18728_/Q _18727_/Q _18726_/Q vssd1 vssd1 vccd1 vccd1 _09153_/D sky130_fd_sc_hd__or3_4
XFILLER_148_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09083_ _09083_/A _17837_/Q _17834_/Q vssd1 vssd1 vccd1 vccd1 _09084_/A sky130_fd_sc_hd__and3_2
XFILLER_175_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09985_ _10089_/S vssd1 vssd1 vccd1 vccd1 _09986_/A sky130_fd_sc_hd__buf_2
XTAP_5107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08936_ _11018_/A vssd1 vssd1 vccd1 vccd1 _08941_/A sky130_fd_sc_hd__buf_12
XTAP_5129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_229_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_8_wb_clk_i clkbuf_5_4_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17939_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_199_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_225_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10760_ _10689_/A _10759_/X _10766_/A vssd1 vssd1 vccd1 vccd1 _10760_/X sky130_fd_sc_hd__a21o_1
XFILLER_213_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09419_ _09419_/A _09419_/B _09419_/C vssd1 vssd1 vccd1 vccd1 _09419_/Y sky130_fd_sc_hd__nand3_2
XFILLER_13_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_213_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_203_wb_clk_i clkbuf_5_6_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18980_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_10691_ _10678_/X _10679_/X _10681_/X _10690_/X vssd1 vssd1 vccd1 vccd1 _10691_/X
+ sky130_fd_sc_hd__a31o_1
X_12430_ _12439_/A _12430_/B _12430_/C vssd1 vssd1 vccd1 vccd1 _12432_/B sky130_fd_sc_hd__nand3_1
XFILLER_40_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_225_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12361_ _12361_/A _12495_/A vssd1 vssd1 vccd1 vccd1 _12387_/A sky130_fd_sc_hd__and2_1
XFILLER_51_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14100_ _18647_/Q _13523_/A _13537_/A _18629_/Q vssd1 vssd1 vccd1 vccd1 _14100_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_166_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19107__78 vssd1 vssd1 vccd1 vccd1 _19107__78/HI _19215_/A sky130_fd_sc_hd__conb_1
XFILLER_4_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11312_ _11368_/A _11312_/B _11997_/A vssd1 vssd1 vccd1 vccd1 _11375_/A sky130_fd_sc_hd__and3_1
X_15080_ _15082_/B _15078_/X _15079_/Y _15066_/X vssd1 vssd1 vccd1 vccd1 _18358_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_180_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12292_ _13418_/C _12292_/B vssd1 vssd1 vccd1 vccd1 _12313_/B sky130_fd_sc_hd__nor2_2
XFILLER_5_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14031_ _18236_/Q _13508_/A _14030_/X _18260_/Q vssd1 vssd1 vccd1 vccd1 _14031_/X
+ sky130_fd_sc_hd__a22o_1
X_11243_ _11243_/A _11243_/B _11245_/B vssd1 vssd1 vccd1 vccd1 _11244_/A sky130_fd_sc_hd__and3_1
XFILLER_106_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11174_ _11177_/B _11198_/B _11174_/C vssd1 vssd1 vccd1 vccd1 _11175_/A sky130_fd_sc_hd__and3b_1
XFILLER_122_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_1178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_164_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10125_ _18127_/Q _10129_/B _10124_/Y vssd1 vssd1 vccd1 vccd1 _10131_/B sky130_fd_sc_hd__a21oi_4
XFILLER_95_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18770_ _18773_/CLK _18770_/D vssd1 vssd1 vccd1 vccd1 _18770_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_67_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15982_ _15982_/A _15993_/B vssd1 vssd1 vccd1 vccd1 _15991_/B sky130_fd_sc_hd__nor2_2
XFILLER_121_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17721_ _17723_/A _19006_/Q vssd1 vssd1 vccd1 vccd1 _17722_/A sky130_fd_sc_hd__and2_1
X_14933_ _14935_/B _14931_/X _14932_/Y _14922_/X vssd1 vssd1 vccd1 vccd1 _18322_/D
+ sky130_fd_sc_hd__o211a_1
X_10056_ _09170_/B _10039_/A _09999_/A _09203_/C vssd1 vssd1 vccd1 vccd1 _10056_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_5674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17652_ _17659_/A _17652_/B vssd1 vssd1 vccd1 vccd1 _17653_/A sky130_fd_sc_hd__and2_1
XFILLER_169_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14864_ _18149_/Q _15015_/B vssd1 vssd1 vccd1 vccd1 _14977_/A sky130_fd_sc_hd__nand2_4
XTAP_4984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16603_ _16621_/A vssd1 vssd1 vccd1 vccd1 _16617_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_223_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13815_ _18924_/Q _13752_/A _13721_/A _18942_/Q vssd1 vssd1 vccd1 vccd1 _13815_/X
+ sky130_fd_sc_hd__a22o_1
X_14795_ _18325_/Q _18289_/Q _14809_/S vssd1 vssd1 vccd1 vccd1 _14795_/X sky130_fd_sc_hd__mux2_1
XFILLER_28_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17583_ _17567_/X _17576_/Y _17582_/X _17577_/Y _18958_/Q vssd1 vssd1 vccd1 vccd1
+ _17584_/B sky130_fd_sc_hd__a32o_1
XFILLER_182_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16534_ _18739_/Q _18703_/Q _16546_/S vssd1 vssd1 vccd1 vccd1 _16534_/X sky130_fd_sc_hd__mux2_1
X_13746_ _18309_/Q _13733_/X _13737_/X _13745_/X vssd1 vssd1 vccd1 vccd1 _13746_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_1_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10958_ _10944_/S _10955_/X _10957_/X _12068_/A vssd1 vssd1 vccd1 vccd1 _10958_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_32_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_231_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_91_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16465_ _16464_/B _16462_/X _16464_/Y _16456_/X vssd1 vssd1 vccd1 vccd1 _18686_/D
+ sky130_fd_sc_hd__o211a_1
X_13677_ _13677_/A vssd1 vssd1 vccd1 vccd1 _13677_/X sky130_fd_sc_hd__buf_6
XFILLER_31_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10889_ _10678_/X _12094_/A _10863_/X _10888_/X _14330_/A vssd1 vssd1 vccd1 vccd1
+ _10889_/X sky130_fd_sc_hd__a311o_1
X_18204_ _18204_/CLK _18204_/D vssd1 vssd1 vccd1 vccd1 _18204_/Q sky130_fd_sc_hd__dfxtp_1
X_15416_ _18473_/Q _18437_/Q _15435_/S vssd1 vssd1 vccd1 vccd1 _15416_/X sky130_fd_sc_hd__mux2_1
X_12628_ _12628_/A _12628_/B vssd1 vssd1 vccd1 vccd1 _12632_/A sky130_fd_sc_hd__nand2_1
X_16396_ _18705_/Q _18669_/Q _16400_/S vssd1 vssd1 vccd1 vccd1 _16396_/X sky130_fd_sc_hd__mux2_1
X_19184_ _19184_/A _09000_/Y vssd1 vssd1 vccd1 vccd1 io_out[22] sky130_fd_sc_hd__ebufn_8
XFILLER_185_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_185_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15347_ _15352_/B _15344_/X _15346_/X _15340_/X vssd1 vssd1 vccd1 vccd1 _18420_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_157_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18135_ _18244_/CLK _18135_/D vssd1 vssd1 vccd1 vccd1 _18135_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_145_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12559_ _12809_/A _12523_/X _12557_/Y _12558_/X _12548_/X vssd1 vssd1 vccd1 vccd1
+ _17919_/D sky130_fd_sc_hd__a221o_1
XFILLER_157_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15278_ _18444_/Q _18408_/Q _15285_/S vssd1 vssd1 vccd1 vccd1 _15278_/X sky130_fd_sc_hd__mux2_1
XFILLER_156_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18066_ _18072_/CLK _18066_/D vssd1 vssd1 vccd1 vccd1 _18066_/Q sky130_fd_sc_hd__dfxtp_1
X_17017_ _18853_/Q _18817_/Q _17026_/S vssd1 vssd1 vccd1 vccd1 _17017_/X sky130_fd_sc_hd__mux2_1
X_14229_ _14283_/A vssd1 vssd1 vccd1 vccd1 _14229_/X sky130_fd_sc_hd__clkbuf_2
Xclkbuf_leaf_78_wb_clk_i clkbuf_5_23_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18633_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_172_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_1302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19121__92 vssd1 vssd1 vccd1 vccd1 _19121__92/HI _19229_/A sky130_fd_sc_hd__conb_1
XFILLER_140_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_112_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09770_ _18107_/Q _10611_/B vssd1 vssd1 vccd1 vccd1 _09785_/B sky130_fd_sc_hd__xnor2_2
XFILLER_100_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18968_ _18980_/CLK _18968_/D vssd1 vssd1 vccd1 vccd1 _18968_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_85_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_140_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17919_ _17919_/CLK _17919_/D vssd1 vssd1 vccd1 vccd1 _17919_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18899_ _18899_/CLK _18899_/D vssd1 vssd1 vccd1 vccd1 _18899_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_66_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_227_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_96_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_226_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_215_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_226_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_208_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_228_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_228_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_224_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_1306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_194_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09204_ _09204_/A _09204_/B _09204_/C vssd1 vssd1 vccd1 vccd1 _09221_/B sky130_fd_sc_hd__nand3_4
XFILLER_22_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_195_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_183_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09135_ _18836_/Q _18835_/Q _18834_/Q vssd1 vssd1 vccd1 vccd1 _09136_/D sky130_fd_sc_hd__or3_4
XFILLER_120_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_202_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09066_ _09066_/A vssd1 vssd1 vccd1 vccd1 _19176_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_147_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_159_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_200_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_1318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_231_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09968_ _09376_/A _09386_/B _09381_/A _09376_/D _12123_/A _14240_/B vssd1 vssd1 vccd1
+ vccd1 _09968_/X sky130_fd_sc_hd__mux4_1
XFILLER_131_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09899_ _10600_/A vssd1 vssd1 vccd1 vccd1 _09972_/B sky130_fd_sc_hd__clkbuf_8
XFILLER_217_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11930_ _11951_/A _11930_/B vssd1 vssd1 vccd1 vccd1 _11979_/A sky130_fd_sc_hd__xnor2_1
XTAP_4269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11861_ _11820_/A _11858_/X _11860_/Y _11852_/X vssd1 vssd1 vccd1 vccd1 _11861_/X
+ sky130_fd_sc_hd__a211o_1
XTAP_2834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13600_ _18729_/Q _13551_/X _13593_/X _13599_/X vssd1 vssd1 vccd1 vccd1 _13600_/X
+ sky130_fd_sc_hd__a211o_1
XTAP_2856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10812_ _09265_/A _09265_/C _10812_/S vssd1 vssd1 vccd1 vccd1 _10812_/X sky130_fd_sc_hd__mux2_1
X_14580_ _16850_/A vssd1 vssd1 vccd1 vccd1 _15184_/A sky130_fd_sc_hd__buf_8
XTAP_2878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11792_ _11790_/X _11791_/X _11789_/Y _11740_/C vssd1 vssd1 vccd1 vccd1 _11792_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_220_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13531_ _13531_/A vssd1 vssd1 vccd1 vccd1 _13532_/A sky130_fd_sc_hd__buf_6
X_10743_ _10743_/A _10743_/B vssd1 vssd1 vccd1 vccd1 _10743_/X sky130_fd_sc_hd__or2_1
XFILLER_198_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_207_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16250_ _18670_/Q _18634_/Q _16250_/S vssd1 vssd1 vccd1 vccd1 _16250_/X sky130_fd_sc_hd__mux2_1
X_13462_ _17840_/Q _13457_/X _13459_/X vssd1 vssd1 vccd1 vccd1 _13463_/B sky130_fd_sc_hd__a21oi_1
XFILLER_174_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10674_ _10706_/B _10705_/A vssd1 vssd1 vccd1 vccd1 _10820_/B sky130_fd_sc_hd__or2b_2
X_15201_ _15250_/A vssd1 vssd1 vccd1 vccd1 _15226_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_16_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12413_ _12414_/A _12414_/B _12414_/C vssd1 vssd1 vccd1 vccd1 _12413_/X sky130_fd_sc_hd__o21a_1
X_16181_ _16181_/A _16773_/B _16181_/C vssd1 vssd1 vccd1 vccd1 _16181_/X sky130_fd_sc_hd__or3_1
X_13393_ _18122_/Q _11021_/X _13337_/X _13383_/X vssd1 vssd1 vccd1 vccd1 _18122_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_182_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15132_ _15182_/A _15132_/B vssd1 vssd1 vccd1 vccd1 _15132_/Y sky130_fd_sc_hd__nand2_1
XFILLER_127_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12344_ _11478_/Y _12336_/X _11473_/Y vssd1 vssd1 vccd1 vccd1 _12346_/B sky130_fd_sc_hd__o21a_1
XFILLER_181_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_177_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15063_ _15527_/A _15136_/C vssd1 vssd1 vccd1 vccd1 _15072_/B sky130_fd_sc_hd__nor2_2
XFILLER_99_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12275_ _11563_/B _12274_/Y _12272_/X vssd1 vssd1 vccd1 vccd1 _17868_/D sky130_fd_sc_hd__o21a_1
X_14014_ _14014_/A vssd1 vssd1 vccd1 vccd1 _14015_/A sky130_fd_sc_hd__clkbuf_8
X_11226_ _17816_/Q _11215_/B _11224_/A _17818_/Q vssd1 vssd1 vccd1 vccd1 _11227_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_4_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_218_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_214_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18822_ _18858_/CLK _18822_/D vssd1 vssd1 vccd1 vccd1 _18822_/Q sky130_fd_sc_hd__dfxtp_2
X_11157_ _17804_/Q vssd1 vssd1 vccd1 vccd1 _11501_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_1_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_209_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10108_ _09711_/A _10093_/X _10107_/X _09657_/X vssd1 vssd1 vccd1 vccd1 _10108_/X
+ sky130_fd_sc_hd__a22o_1
X_18753_ _18788_/CLK _18753_/D vssd1 vssd1 vccd1 vccd1 _18753_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_95_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15965_ _15971_/B _15963_/X _15964_/X _15948_/X vssd1 vssd1 vccd1 vccd1 _18567_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_5460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11088_ _11088_/A vssd1 vssd1 vccd1 vccd1 _17791_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_62_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17704_ _17704_/A _17704_/B vssd1 vssd1 vccd1 vccd1 _17704_/Y sky130_fd_sc_hd__nor2_1
XFILLER_209_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14916_ _16431_/A vssd1 vssd1 vccd1 vccd1 _15527_/A sky130_fd_sc_hd__buf_4
X_10039_ _10039_/A vssd1 vssd1 vccd1 vccd1 _10040_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_3_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18684_ _18686_/CLK _18684_/D vssd1 vssd1 vccd1 vccd1 _18684_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_63_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_196_wb_clk_i _18176_/CLK vssd1 vssd1 vccd1 vccd1 _19000_/CLK sky130_fd_sc_hd__clkbuf_16
X_15896_ _18589_/Q _18553_/Q _15899_/S vssd1 vssd1 vccd1 vccd1 _15896_/X sky130_fd_sc_hd__mux2_1
XTAP_4770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17635_ _17635_/A _17663_/B vssd1 vssd1 vccd1 vccd1 _17635_/Y sky130_fd_sc_hd__nor2_1
XFILLER_75_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_125_wb_clk_i clkbuf_5_25_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18416_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_184_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14847_ _14849_/B _14845_/X _14846_/Y _14839_/X vssd1 vssd1 vccd1 vccd1 _18301_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_91_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_223_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17566_ _17640_/A vssd1 vssd1 vccd1 vccd1 _17587_/A sky130_fd_sc_hd__clkbuf_1
X_14778_ _14778_/A vssd1 vssd1 vccd1 vccd1 _14778_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_63_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_223_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_225_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_205_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_5_25_0_wb_clk_i clkbuf_5_25_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_5_25_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_2
X_16517_ _16650_/B vssd1 vssd1 vccd1 vccd1 _16568_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_147_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13729_ _18264_/Q _13714_/X _13698_/A _18255_/Q _13728_/X vssd1 vssd1 vccd1 vccd1
+ _13729_/X sky130_fd_sc_hd__a221o_1
XFILLER_32_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17497_ _17497_/A vssd1 vssd1 vccd1 vccd1 _17497_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_176_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_225_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19236_ _19236_/A _08946_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[36] sky130_fd_sc_hd__ebufn_8
XFILLER_56_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16448_ _16450_/B _16446_/X _16447_/Y _16437_/X vssd1 vssd1 vccd1 vccd1 _18682_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_165_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19167_ _19167_/A _09031_/Y vssd1 vssd1 vccd1 vccd1 io_out[5] sky130_fd_sc_hd__ebufn_8
X_16379_ _18665_/Q _16378_/B _16378_/Y _16376_/X vssd1 vssd1 vccd1 vccd1 _18665_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_219_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18118_ _18125_/CLK _18118_/D vssd1 vssd1 vccd1 vccd1 _18118_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_173_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18049_ _18072_/CLK _18049_/D vssd1 vssd1 vccd1 vccd1 _18049_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_145_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19098__69 vssd1 vssd1 vccd1 vccd1 _19098__69/HI _19206_/A sky130_fd_sc_hd__conb_1
XFILLER_132_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09822_ _09822_/A _09844_/A vssd1 vssd1 vccd1 vccd1 _09843_/A sky130_fd_sc_hd__nand2_1
XFILLER_8_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_150_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_230_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09753_ _09753_/A _09753_/B vssd1 vssd1 vccd1 vccd1 _09764_/A sky130_fd_sc_hd__nand2_1
XFILLER_104_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09684_ _09684_/A _09684_/B vssd1 vssd1 vccd1 vccd1 _09704_/B sky130_fd_sc_hd__and2_1
XFILLER_227_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_211_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_195_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_168_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09118_ _18767_/Q _18766_/Q _18765_/Q vssd1 vssd1 vccd1 vccd1 _10350_/A sky130_fd_sc_hd__or3_4
XFILLER_129_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10390_ _09354_/C _09971_/S _10389_/X _09937_/X vssd1 vssd1 vccd1 vccd1 _10390_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_164_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09049_ _09052_/A vssd1 vssd1 vccd1 vccd1 _09049_/Y sky130_fd_sc_hd__inv_2
XFILLER_159_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12060_ _09683_/X _13526_/B _12058_/X _12059_/Y vssd1 vssd1 vccd1 vccd1 _12060_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_104_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11011_ _17814_/Q _11190_/A _11011_/C _11011_/D vssd1 vssd1 vccd1 vccd1 _11012_/A
+ sky130_fd_sc_hd__or4_1
XFILLER_77_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_219_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_219_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15750_ _18553_/Q _18517_/Q _15753_/S vssd1 vssd1 vccd1 vccd1 _15750_/X sky130_fd_sc_hd__mux2_1
XTAP_4055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12962_ _12962_/A _12969_/B vssd1 vssd1 vccd1 vccd1 _12962_/Y sky130_fd_sc_hd__nor2_1
XTAP_4066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_50 _10541_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_61 _17747_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_72 _13532_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_83 _13596_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14701_ _18266_/Q _14700_/B _14700_/Y _14692_/X vssd1 vssd1 vccd1 vccd1 _18266_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_3343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11913_ _10256_/A _18128_/Q _11913_/S vssd1 vssd1 vccd1 vccd1 _11913_/X sky130_fd_sc_hd__mux2_1
XTAP_4099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15681_ _15720_/A vssd1 vssd1 vccd1 vccd1 _15681_/X sky130_fd_sc_hd__clkbuf_2
XINSDIODE2_94 _14124_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12893_ _12792_/X _12895_/C _12874_/X vssd1 vssd1 vccd1 vccd1 _12893_/Y sky130_fd_sc_hd__o21ai_1
XTAP_2620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17420_ _17420_/A vssd1 vssd1 vccd1 vccd1 _17497_/A sky130_fd_sc_hd__clkbuf_2
XTAP_2653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14632_ _14681_/A _14635_/B vssd1 vssd1 vccd1 vccd1 _14632_/Y sky130_fd_sc_hd__nand2_1
XTAP_3398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11844_ _11844_/A _11844_/B _11842_/A vssd1 vssd1 vccd1 vccd1 _11845_/C sky130_fd_sc_hd__or3b_1
XFILLER_92_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14563_ _18174_/Q _18173_/Q _18169_/Q _18170_/Q vssd1 vssd1 vccd1 vccd1 _14672_/A
+ sky130_fd_sc_hd__or4b_2
X_17351_ _17491_/A _17351_/B vssd1 vssd1 vccd1 vccd1 _17360_/B sky130_fd_sc_hd__nor2_2
X_11775_ _11775_/A vssd1 vssd1 vccd1 vccd1 _11781_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_220_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16302_ _16325_/A _16305_/B vssd1 vssd1 vccd1 vccd1 _16302_/Y sky130_fd_sc_hd__nand2_1
XTAP_1996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13514_ _13582_/A vssd1 vssd1 vccd1 vccd1 _13515_/A sky130_fd_sc_hd__buf_4
X_10726_ _09114_/B _09109_/B _09119_/C _09109_/C _10695_/A _10764_/A vssd1 vssd1 vccd1
+ vccd1 _10726_/X sky130_fd_sc_hd__mux4_2
XFILLER_207_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14494_ _18221_/Q _14502_/B vssd1 vssd1 vccd1 vccd1 _14495_/A sky130_fd_sc_hd__and2_1
XFILLER_9_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17282_ _17318_/A _17425_/B _17318_/C vssd1 vssd1 vccd1 vccd1 _17282_/X sky130_fd_sc_hd__or3_1
XFILLER_140_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19021_ _19021_/CLK _19021_/D vssd1 vssd1 vccd1 vccd1 _19021_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_174_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16233_ _18140_/Q _16528_/B vssd1 vssd1 vccd1 vccd1 _16348_/A sky130_fd_sc_hd__nand2_1
X_13445_ _13441_/X _13443_/Y _13444_/X _13428_/Y vssd1 vssd1 vccd1 vccd1 _13455_/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_16_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10657_ _10721_/A vssd1 vssd1 vccd1 vccd1 _10813_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_167_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16164_ _16919_/A vssd1 vssd1 vccd1 vccd1 _16757_/A sky130_fd_sc_hd__buf_6
XFILLER_155_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13376_ _13346_/X _13374_/Y _13379_/B vssd1 vssd1 vccd1 vccd1 _18110_/D sky130_fd_sc_hd__a21boi_1
XFILLER_186_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10588_ _10009_/A _10586_/X _10587_/X _10040_/A vssd1 vssd1 vccd1 vccd1 _10588_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_155_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15115_ _15115_/A _15118_/B vssd1 vssd1 vccd1 vccd1 _15115_/Y sky130_fd_sc_hd__nand2_1
XFILLER_154_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12327_ _12327_/A _12327_/B _12327_/C vssd1 vssd1 vccd1 vccd1 _12328_/B sky130_fd_sc_hd__and3_1
XFILLER_86_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16095_ _18635_/Q _18599_/Q _16113_/S vssd1 vssd1 vccd1 vccd1 _16095_/X sky130_fd_sc_hd__mux2_1
XFILLER_170_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15046_ _15083_/A vssd1 vssd1 vccd1 vccd1 _15046_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_141_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12258_ _17864_/Q _13066_/B _12258_/C vssd1 vssd1 vccd1 vccd1 _12259_/A sky130_fd_sc_hd__and3_1
XFILLER_107_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_1335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_218_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11209_ _11209_/A _11209_/B vssd1 vssd1 vccd1 vccd1 _11210_/C sky130_fd_sc_hd__or2_1
XFILLER_122_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12189_ _12470_/B vssd1 vssd1 vccd1 vccd1 _12499_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_214_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_229_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18805_ _18806_/CLK _18805_/D vssd1 vssd1 vccd1 vccd1 _18805_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_110_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16997_ _18848_/Q _18812_/Q _17005_/S vssd1 vssd1 vccd1 vccd1 _16997_/X sky130_fd_sc_hd__mux2_1
XFILLER_23_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18736_ _18765_/CLK _18736_/D vssd1 vssd1 vccd1 vccd1 _18736_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_97_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15948_ _16028_/A vssd1 vssd1 vccd1 vccd1 _15948_/X sky130_fd_sc_hd__clkbuf_2
XTAP_5290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_224_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_225_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18667_ _18683_/CLK _18667_/D vssd1 vssd1 vccd1 vccd1 _18667_/Q sky130_fd_sc_hd__dfxtp_2
X_15879_ _18585_/Q _18549_/Q _15879_/S vssd1 vssd1 vccd1 vccd1 _15879_/X sky130_fd_sc_hd__mux2_1
XFILLER_97_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17618_ _14354_/X _14612_/X _17547_/X _17617_/X _17556_/X vssd1 vssd1 vccd1 vccd1
+ _18966_/D sky130_fd_sc_hd__o311a_1
XFILLER_197_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18598_ _18608_/CLK _18598_/D vssd1 vssd1 vccd1 vccd1 _18598_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_145_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_224_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_225_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17549_ _17549_/A _17549_/B vssd1 vssd1 vccd1 vccd1 _17581_/A sky130_fd_sc_hd__nor2_1
XFILLER_20_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_189_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_1339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_225_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19219_ _19219_/A _08959_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[19] sky130_fd_sc_hd__ebufn_8
XFILLER_177_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_93_wb_clk_i _18144_/CLK vssd1 vssd1 vccd1 vccd1 _18147_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_149_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_22_wb_clk_i clkbuf_5_6_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18908_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_173_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_195_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_219_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09805_ _09805_/A _09805_/B vssd1 vssd1 vccd1 vccd1 _09806_/B sky130_fd_sc_hd__xnor2_1
XFILLER_140_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09736_ _09743_/A _10116_/B _09735_/Y vssd1 vssd1 vccd1 vccd1 _09739_/A sky130_fd_sc_hd__a21bo_1
XFILLER_227_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09667_ _12072_/B _09667_/B vssd1 vssd1 vccd1 vccd1 _09668_/B sky130_fd_sc_hd__xnor2_2
XFILLER_28_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09598_ _09586_/A _09586_/B _09598_/S vssd1 vssd1 vccd1 vccd1 _09610_/A sky130_fd_sc_hd__mux2_2
XFILLER_91_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_230_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_231_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_208_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11560_ _11622_/A _11554_/X _11559_/X vssd1 vssd1 vccd1 vccd1 _11560_/X sky130_fd_sc_hd__a21o_1
XFILLER_11_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10511_ _09098_/D _09103_/C _09103_/A _09093_/D _10464_/X _10235_/A vssd1 vssd1 vccd1
+ vccd1 _10512_/C sky130_fd_sc_hd__mux4_2
XFILLER_10_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11491_ _11491_/A vssd1 vssd1 vccd1 vccd1 _11491_/Y sky130_fd_sc_hd__inv_2
XFILLER_7_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_196_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13230_ _13230_/A vssd1 vssd1 vccd1 vccd1 _18069_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_10_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_196_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_1302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10442_ _12031_/A _14289_/A vssd1 vssd1 vccd1 vccd1 _10443_/A sky130_fd_sc_hd__and2_4
XFILLER_108_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13161_ _13161_/A vssd1 vssd1 vccd1 vccd1 _18038_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_13_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_1305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10373_ _09337_/A _09332_/C _09327_/D _09337_/D _09953_/A _10349_/S vssd1 vssd1 vccd1
+ vccd1 _10374_/B sky130_fd_sc_hd__mux4_1
XFILLER_87_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12112_ _12112_/A _12112_/B _12112_/C vssd1 vssd1 vccd1 vccd1 _12112_/X sky130_fd_sc_hd__and3_1
XFILLER_174_1338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13092_ _18007_/Q _14377_/A vssd1 vssd1 vccd1 vccd1 _13093_/A sky130_fd_sc_hd__or2_1
XFILLER_215_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16920_ _17503_/A _16960_/B vssd1 vssd1 vccd1 vccd1 _16930_/B sky130_fd_sc_hd__nor2_2
XFILLER_3_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12043_ _12043_/A _12043_/B vssd1 vssd1 vccd1 vccd1 _13693_/A sky130_fd_sc_hd__and2_2
XFILLER_105_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_215_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16851_ _17446_/A _16906_/B vssd1 vssd1 vccd1 vccd1 _16860_/B sky130_fd_sc_hd__nor2_2
XFILLER_131_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15802_ _15815_/A _15806_/B vssd1 vssd1 vccd1 vccd1 _15802_/Y sky130_fd_sc_hd__nand2_1
XFILLER_150_1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16782_ _16779_/B _16778_/X _16779_/Y _16781_/X vssd1 vssd1 vccd1 vccd1 _18764_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_20_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13994_ _18571_/Q _13772_/X _13752_/X _18565_/Q _13993_/X vssd1 vssd1 vccd1 vccd1
+ _13994_/X sky130_fd_sc_hd__a221o_1
XFILLER_46_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18521_ _18546_/CLK _18521_/D vssd1 vssd1 vccd1 vccd1 _18521_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_18_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15733_ _18549_/Q _18513_/Q _15733_/S vssd1 vssd1 vccd1 vccd1 _15733_/X sky130_fd_sc_hd__mux2_1
XFILLER_20_1238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12945_ _12945_/A vssd1 vssd1 vccd1 vccd1 _17972_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_80_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18452_ _18467_/CLK _18452_/D vssd1 vssd1 vccd1 vccd1 _18452_/Q sky130_fd_sc_hd__dfxtp_4
XTAP_3184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15664_ _15962_/A _15696_/B vssd1 vssd1 vccd1 vccd1 _15673_/B sky130_fd_sc_hd__nor2_1
XFILLER_206_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12876_ _12824_/A _12877_/C _12875_/Y vssd1 vssd1 vccd1 vccd1 _17955_/D sky130_fd_sc_hd__a21oi_1
XTAP_2461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17403_ _17464_/A vssd1 vssd1 vccd1 vccd1 _17453_/A sky130_fd_sc_hd__clkbuf_2
X_14615_ _14608_/X _14612_/A _18247_/Q vssd1 vssd1 vccd1 vccd1 _14615_/Y sky130_fd_sc_hd__o21bai_1
XTAP_2483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18383_ _18392_/CLK _18383_/D vssd1 vssd1 vccd1 vccd1 _18383_/Q sky130_fd_sc_hd__dfxtp_2
X_11827_ _11778_/X _11825_/Y _11826_/X _11809_/X vssd1 vssd1 vccd1 vccd1 _11827_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_57_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15595_ _15616_/A vssd1 vssd1 vccd1 vccd1 _15595_/X sky130_fd_sc_hd__clkbuf_2
XTAP_1760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17334_ _17334_/A _17336_/B vssd1 vssd1 vccd1 vccd1 _17334_/Y sky130_fd_sc_hd__nand2_1
XFILLER_222_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14546_ _18233_/Q _14545_/B _14545_/Y _14533_/X vssd1 vssd1 vccd1 vccd1 _18233_/D
+ sky130_fd_sc_hd__o211a_1
X_11758_ _11729_/X _11730_/Y _11752_/X _11757_/Y vssd1 vssd1 vccd1 vccd1 _11758_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_81_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_230_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_187_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10709_ _10622_/Y _10673_/X _10910_/C _10691_/X _10708_/X vssd1 vssd1 vccd1 vccd1
+ _10709_/X sky130_fd_sc_hd__a221o_1
XFILLER_31_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17265_ _17265_/A _17549_/B vssd1 vssd1 vccd1 vccd1 _17331_/A sky130_fd_sc_hd__or2_1
XFILLER_105_1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11689_ _11689_/A _11700_/A vssd1 vssd1 vccd1 vccd1 _11689_/Y sky130_fd_sc_hd__nand2_1
X_14477_ _14477_/A vssd1 vssd1 vccd1 vccd1 _18213_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_179_1216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19004_ _19004_/CLK _19004_/D vssd1 vssd1 vccd1 vccd1 _19004_/Q sky130_fd_sc_hd__dfxtp_1
X_16216_ _16216_/A vssd1 vssd1 vccd1 vccd1 _16268_/A sky130_fd_sc_hd__buf_2
X_13428_ _11070_/X _13422_/Y _13426_/Y _13447_/B vssd1 vssd1 vccd1 vccd1 _13428_/Y
+ sky130_fd_sc_hd__o211ai_2
XFILLER_31_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17196_ _17210_/A _17200_/B vssd1 vssd1 vccd1 vccd1 _17196_/Y sky130_fd_sc_hd__nand2_1
XFILLER_6_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16147_ _16202_/A _16147_/B vssd1 vssd1 vccd1 vccd1 _16147_/Y sky130_fd_sc_hd__nand2_1
XFILLER_155_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13359_ _17778_/Q _17704_/A _13356_/B _12217_/A vssd1 vssd1 vccd1 vccd1 _13363_/B
+ sky130_fd_sc_hd__o31a_1
XFILLER_142_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16078_ _16130_/A _16082_/B vssd1 vssd1 vccd1 vccd1 _16078_/Y sky130_fd_sc_hd__nand2_1
X_19068__39 vssd1 vssd1 vccd1 vccd1 _19068__39/HI _19162_/A sky130_fd_sc_hd__conb_1
XFILLER_143_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15029_ _15172_/A _15085_/B vssd1 vssd1 vccd1 vccd1 _15038_/B sky130_fd_sc_hd__nor2_2
XFILLER_142_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_229_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_140_wb_clk_i clkbuf_5_26_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18324_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_29_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_1299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput2 io_in[10] vssd1 vssd1 vccd1 vccd1 input2/X sky130_fd_sc_hd__buf_8
XFILLER_7_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_216_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09521_ _14319_/S vssd1 vssd1 vccd1 vccd1 _14332_/S sky130_fd_sc_hd__clkbuf_2
X_18719_ _18719_/CLK _18719_/D vssd1 vssd1 vccd1 vccd1 _18719_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_225_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_213_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09452_ _09221_/B _09451_/X _09188_/X vssd1 vssd1 vccd1 vccd1 _09452_/X sky130_fd_sc_hd__a21o_1
XFILLER_52_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_224_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_212_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09383_ _18392_/Q _18391_/Q _18390_/Q vssd1 vssd1 vccd1 vccd1 _09386_/B sky130_fd_sc_hd__or3_4
XFILLER_52_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_165_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_228_wb_clk_i _17864_/CLK vssd1 vssd1 vccd1 vccd1 _17861_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_69_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_1366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19082__53 vssd1 vssd1 vccd1 vccd1 _19082__53/HI _19190_/A sky130_fd_sc_hd__conb_1
XFILLER_101_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09719_ _10582_/S _09719_/B vssd1 vssd1 vccd1 vccd1 _09720_/A sky130_fd_sc_hd__nor2_4
X_10991_ _18997_/Q _10990_/X _10982_/X hold3/X vssd1 vssd1 vccd1 vccd1 _18997_/D sky130_fd_sc_hd__a22o_1
XFILLER_90_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_216_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12730_ _12921_/A vssd1 vssd1 vccd1 vccd1 _12919_/B sky130_fd_sc_hd__clkbuf_2
XTAP_1001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_4_6_0_wb_clk_i clkbuf_4_7_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_4_6_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_231_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12661_ _12662_/A _12662_/B vssd1 vssd1 vccd1 vccd1 _12663_/A sky130_fd_sc_hd__and2_1
XTAP_1056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_231_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_208_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11612_ _17856_/Q vssd1 vssd1 vccd1 vccd1 _11614_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_14400_ _17591_/A _14423_/A vssd1 vssd1 vccd1 vccd1 _14428_/A sky130_fd_sc_hd__or2_1
XFILLER_187_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15380_ _16889_/A vssd1 vssd1 vccd1 vccd1 _15984_/B sky130_fd_sc_hd__buf_2
X_12592_ _12590_/A _12590_/B _12591_/X vssd1 vssd1 vccd1 vccd1 _12592_/X sky130_fd_sc_hd__o21a_1
XFILLER_23_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_230_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_212_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14331_ _14317_/A _12056_/A _14205_/A _10939_/A _14330_/Y vssd1 vssd1 vccd1 vccd1
+ _14331_/X sky130_fd_sc_hd__a221o_1
X_11543_ _13518_/A vssd1 vssd1 vccd1 vccd1 _13526_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_51_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_195_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17050_ _17072_/A _17483_/B _17085_/C vssd1 vssd1 vccd1 vccd1 _17050_/X sky130_fd_sc_hd__or3_1
X_14262_ _14219_/X _14257_/Y _14261_/X _14222_/Y vssd1 vssd1 vccd1 vccd1 _14262_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_156_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11474_ _11459_/A _11478_/B _12340_/A _11473_/Y vssd1 vssd1 vccd1 vccd1 _11474_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_184_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16001_ _16003_/B _15999_/X _16000_/Y _15988_/X vssd1 vssd1 vccd1 vccd1 _18577_/D
+ sky130_fd_sc_hd__o211a_1
X_13213_ _13257_/A vssd1 vssd1 vccd1 vccd1 _13222_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_87_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10425_ _12047_/A vssd1 vssd1 vccd1 vccd1 _10939_/C sky130_fd_sc_hd__buf_2
X_14193_ _18222_/Q _18221_/Q _18220_/Q _18219_/Q vssd1 vssd1 vccd1 vccd1 _14196_/A
+ sky130_fd_sc_hd__or4_1
XFILLER_174_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13144_ _13144_/A vssd1 vssd1 vccd1 vccd1 _18030_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_152_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10356_ _10356_/A _10356_/B vssd1 vssd1 vccd1 vccd1 _10356_/X sky130_fd_sc_hd__or2_1
XFILLER_48_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_1266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13075_ _18001_/Q _12718_/X _13072_/X _13074_/X vssd1 vssd1 vccd1 vccd1 _18001_/D
+ sky130_fd_sc_hd__o211a_1
X_17952_ _17954_/CLK _17952_/D vssd1 vssd1 vccd1 vccd1 _17952_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_111_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_215_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10287_ _09916_/X _10285_/X _10286_/X _09895_/X _09969_/X vssd1 vssd1 vccd1 vccd1
+ _10288_/B sky130_fd_sc_hd__a221o_1
XFILLER_78_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16903_ _16957_/A _16903_/B vssd1 vssd1 vccd1 vccd1 _16903_/Y sky130_fd_sc_hd__nand2_1
X_12026_ _11984_/C _12026_/B _12026_/C _12026_/D vssd1 vssd1 vccd1 vccd1 _12027_/D
+ sky130_fd_sc_hd__and4b_4
X_17883_ _17883_/CLK _17883_/D vssd1 vssd1 vccd1 vccd1 _17883_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_120_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16834_ _16833_/B _16831_/X _16833_/Y _16825_/X vssd1 vssd1 vccd1 vccd1 _18776_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_120_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_219_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16765_ _16769_/B _16762_/X _16764_/Y _16760_/X vssd1 vssd1 vccd1 vccd1 _18760_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_18_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13977_ _18301_/Q _13759_/X _13780_/X _18292_/Q _13976_/X vssd1 vssd1 vccd1 vccd1
+ _13977_/X sky130_fd_sc_hd__a221o_4
XFILLER_20_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18504_ _18504_/CLK _18504_/D vssd1 vssd1 vccd1 vccd1 _18504_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_46_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15716_ _15719_/B _15714_/X _15715_/Y _15700_/X vssd1 vssd1 vccd1 vccd1 _18508_/D
+ sky130_fd_sc_hd__o211a_1
X_12928_ _12748_/A _12924_/Y _12927_/Y vssd1 vssd1 vccd1 vccd1 _12928_/X sky130_fd_sc_hd__o21a_1
XFILLER_59_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16696_ _16699_/B _16694_/X _16695_/Y _16683_/X vssd1 vssd1 vccd1 vccd1 _18742_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_34_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18435_ _18443_/CLK _18435_/D vssd1 vssd1 vccd1 vccd1 _18435_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_22_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_221_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15647_ _15717_/A vssd1 vssd1 vccd1 vccd1 _15665_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_185_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_222_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12859_ _12865_/C _12859_/B _12874_/A vssd1 vssd1 vccd1 vccd1 _12860_/A sky130_fd_sc_hd__and3b_1
XTAP_2291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18366_ _18380_/CLK _18366_/D vssd1 vssd1 vccd1 vccd1 _18366_/Q sky130_fd_sc_hd__dfxtp_2
X_15578_ _15578_/A vssd1 vssd1 vccd1 vccd1 _15630_/A sky130_fd_sc_hd__clkbuf_2
XTAP_1590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17317_ _18927_/Q _18891_/Q _17317_/S vssd1 vssd1 vccd1 vccd1 _17317_/X sky130_fd_sc_hd__mux2_1
XFILLER_186_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14529_ _14702_/A vssd1 vssd1 vccd1 vccd1 _17412_/A sky130_fd_sc_hd__buf_4
X_18297_ _18308_/CLK _18297_/D vssd1 vssd1 vccd1 vccd1 _18297_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_147_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17248_ _18910_/Q _18874_/Q _17262_/S vssd1 vssd1 vccd1 vccd1 _17248_/X sky130_fd_sc_hd__mux2_1
XFILLER_174_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17179_ _18893_/Q _18857_/Q _17199_/S vssd1 vssd1 vccd1 vccd1 _17179_/X sky130_fd_sc_hd__mux2_1
XFILLER_227_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_1322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08952_ _08954_/A vssd1 vssd1 vccd1 vccd1 _08952_/Y sky130_fd_sc_hd__inv_2
XFILLER_131_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09504_ _18203_/Q _18202_/Q _14445_/B vssd1 vssd1 vccd1 vccd1 _09505_/B sky130_fd_sc_hd__or3_1
XFILLER_53_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_213_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_213_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09435_ _09435_/A _09435_/B vssd1 vssd1 vccd1 vccd1 _09475_/A sky130_fd_sc_hd__nor2_1
XFILLER_38_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_212_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_205_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09366_ _18284_/Q _18283_/Q _18282_/Q vssd1 vssd1 vccd1 vccd1 _09370_/A sky130_fd_sc_hd__or3_2
XFILLER_200_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_200_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_205_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09297_ _18488_/Q _18487_/Q _18486_/Q vssd1 vssd1 vccd1 vccd1 _09299_/C sky130_fd_sc_hd__or3_2
XFILLER_165_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_166_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_opt_1_0_wb_clk_i _18254_/CLK vssd1 vssd1 vccd1 vccd1 clkbuf_opt_1_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_84_1305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10210_ _10210_/A _10210_/B vssd1 vssd1 vccd1 vccd1 _10211_/B sky130_fd_sc_hd__and2_1
XFILLER_134_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_97_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11190_ _11190_/A _11196_/D vssd1 vssd1 vccd1 vccd1 _11193_/B sky130_fd_sc_hd__nand2_1
XFILLER_161_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10141_ _10141_/A _10141_/B vssd1 vssd1 vccd1 vccd1 _10144_/A sky130_fd_sc_hd__xnor2_2
XFILLER_106_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10072_ _09227_/A _09237_/B _10826_/A _09227_/D _10004_/B _10025_/X vssd1 vssd1 vccd1
+ vccd1 _10072_/X sky130_fd_sc_hd__mux4_1
XTAP_5834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13900_ _18553_/Q _13906_/B vssd1 vssd1 vccd1 vccd1 _13900_/X sky130_fd_sc_hd__and2_1
XTAP_5867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14880_ _14919_/A _15175_/B _14906_/C vssd1 vssd1 vccd1 vccd1 _14880_/X sky130_fd_sc_hd__or3_1
XTAP_5889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_229_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13831_ _13572_/X _13610_/X _13830_/X _18166_/Q _14222_/A vssd1 vssd1 vccd1 vccd1
+ _13832_/B sky130_fd_sc_hd__o32a_2
XFILLER_46_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16550_ _18743_/Q _18707_/Q _16565_/S vssd1 vssd1 vccd1 vccd1 _16550_/X sky130_fd_sc_hd__mux2_1
XINSDIODE2_208 _13531_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13762_ _18498_/Q _13715_/X _13734_/X _18492_/Q _13761_/X vssd1 vssd1 vccd1 vccd1
+ _13762_/X sky130_fd_sc_hd__a221o_1
XFILLER_28_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10974_ _13415_/A _13415_/B _13412_/C _13418_/B vssd1 vssd1 vccd1 vccd1 _14282_/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_16_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINSDIODE2_219 _13780_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15501_ _15500_/B _15499_/X _15500_/Y _15496_/X vssd1 vssd1 vccd1 vccd1 _18455_/D
+ sky130_fd_sc_hd__o211a_1
XPHY_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12713_ _14185_/A _12713_/B vssd1 vssd1 vccd1 vccd1 _17939_/D sky130_fd_sc_hd__nand2_1
XFILLER_203_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16481_ _16491_/A _16773_/B _16481_/C vssd1 vssd1 vccd1 vccd1 _16481_/X sky130_fd_sc_hd__or3_1
XFILLER_204_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13693_ _13693_/A _13710_/C vssd1 vssd1 vccd1 vccd1 _13693_/Y sky130_fd_sc_hd__nor2_8
X_18220_ _18222_/CLK _18220_/D vssd1 vssd1 vccd1 vccd1 _18220_/Q sky130_fd_sc_hd__dfxtp_1
X_15432_ _15431_/B _15430_/X _15431_/Y _15428_/X vssd1 vssd1 vccd1 vccd1 _18440_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_62_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12644_ _17932_/Q vssd1 vssd1 vccd1 vccd1 _12646_/A sky130_fd_sc_hd__clkinv_2
XFILLER_197_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18151_ _18151_/CLK _18151_/D vssd1 vssd1 vccd1 vccd1 _18151_/Q sky130_fd_sc_hd__dfxtp_1
X_15363_ _15404_/A vssd1 vssd1 vccd1 vccd1 _15363_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_12575_ _12575_/A _12575_/B vssd1 vssd1 vccd1 vccd1 _12575_/Y sky130_fd_sc_hd__nor2_1
XFILLER_129_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17102_ _17105_/B _17099_/X _17101_/Y _17096_/X vssd1 vssd1 vccd1 vccd1 _18838_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_200_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14314_ _18177_/Q vssd1 vssd1 vccd1 vccd1 _15903_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_89_1216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11526_ _11701_/A _11526_/B _11512_/C vssd1 vssd1 vccd1 vccd1 _11526_/X sky130_fd_sc_hd__or3b_1
X_18082_ _18087_/CLK _18082_/D vssd1 vssd1 vccd1 vccd1 _18082_/Q sky130_fd_sc_hd__dfxtp_1
X_15294_ _16566_/A vssd1 vssd1 vccd1 vccd1 _15562_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_102_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17033_ _17035_/B _17031_/X _17032_/Y _17020_/X vssd1 vssd1 vccd1 vccd1 _18820_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_172_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11457_ _17886_/Q vssd1 vssd1 vccd1 vccd1 _11479_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_14245_ _14243_/X _14227_/X _14229_/X _14244_/X _18170_/Q vssd1 vssd1 vccd1 vccd1
+ _14245_/X sky130_fd_sc_hd__a311o_1
XFILLER_171_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10408_ _10513_/A vssd1 vssd1 vccd1 vccd1 _10936_/S sky130_fd_sc_hd__clkbuf_2
X_14176_ _18677_/Q _13492_/A _13500_/A _18692_/Q vssd1 vssd1 vccd1 vccd1 _14176_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_194_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11388_ _11388_/A _11388_/B vssd1 vssd1 vccd1 vccd1 _11388_/Y sky130_fd_sc_hd__nor2_1
XFILLER_152_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10339_ _09114_/B _09109_/B _09119_/C _09109_/C _10286_/S _14240_/B vssd1 vssd1 vccd1
+ vccd1 _10339_/X sky130_fd_sc_hd__mux4_1
XFILLER_124_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13127_ _13129_/A _18024_/Q vssd1 vssd1 vccd1 vccd1 _13128_/A sky130_fd_sc_hd__and2_1
XFILLER_113_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18984_ _18986_/CLK _18984_/D vssd1 vssd1 vccd1 vccd1 _18984_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_97_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13058_ _13054_/Y _13058_/B vssd1 vssd1 vccd1 vccd1 _13063_/A sky130_fd_sc_hd__and2b_1
X_17935_ _17939_/CLK _17935_/D vssd1 vssd1 vccd1 vccd1 _17935_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_87_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12009_ _12048_/A _13421_/A _12009_/C _12009_/D vssd1 vssd1 vccd1 vccd1 _12010_/D
+ sky130_fd_sc_hd__and4b_1
XFILLER_113_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17866_ _19032_/CLK _17866_/D vssd1 vssd1 vccd1 vccd1 _17866_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_94_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16817_ _16817_/A vssd1 vssd1 vccd1 vccd1 _17423_/A sky130_fd_sc_hd__buf_4
XFILLER_213_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17797_ _17851_/CLK _17797_/D vssd1 vssd1 vccd1 vccd1 _17797_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_19_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16748_ _16808_/A vssd1 vssd1 vccd1 vccd1 _16796_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_19_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16679_ _16686_/B _16677_/X _16678_/X _16659_/X vssd1 vssd1 vccd1 vccd1 _18738_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_61_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09220_ _09220_/A _09220_/B _09220_/C vssd1 vssd1 vccd1 vccd1 _09430_/D sky130_fd_sc_hd__nand3_1
XFILLER_22_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18418_ _18423_/CLK _18418_/D vssd1 vssd1 vccd1 vccd1 _18418_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_107_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_226_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09151_ _18701_/Q _18700_/Q _18699_/Q vssd1 vssd1 vccd1 vccd1 _10722_/A sky130_fd_sc_hd__or3_4
X_18349_ _18356_/CLK _18349_/D vssd1 vssd1 vccd1 vccd1 _18349_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_147_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09082_ _09082_/A vssd1 vssd1 vccd1 vccd1 _19179_/A sky130_fd_sc_hd__buf_2
XFILLER_174_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_190_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_190_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_162_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_200_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09984_ _10060_/A vssd1 vssd1 vccd1 vccd1 _10089_/S sky130_fd_sc_hd__buf_6
XFILLER_104_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08935_ _08935_/A vssd1 vssd1 vccd1 vccd1 _08935_/Y sky130_fd_sc_hd__inv_2
XFILLER_76_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_69_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_1363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_229_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19052__23 vssd1 vssd1 vccd1 vccd1 _19052__23/HI _19146_/A sky130_fd_sc_hd__conb_1
XTAP_3739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_198_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_213_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_1292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09418_ _09418_/A _09418_/B _09418_/C _09418_/D vssd1 vssd1 vccd1 vccd1 _09419_/C
+ sky130_fd_sc_hd__and4_1
XFILLER_201_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10690_ _10864_/A _10679_/A _10684_/X _10689_/X vssd1 vssd1 vccd1 vccd1 _10690_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_13_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_1208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09349_ _09349_/A _09349_/B _10391_/A _09349_/D vssd1 vssd1 vccd1 vccd1 _09355_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_40_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_205_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12360_ _12147_/X _12353_/Y _12495_/A _12359_/X vssd1 vssd1 vccd1 vccd1 _17892_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_32_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_218_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11311_ _11970_/C _11806_/B vssd1 vssd1 vccd1 vccd1 _11997_/A sky130_fd_sc_hd__nor2_2
XFILLER_126_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12291_ _12327_/A vssd1 vssd1 vccd1 vccd1 _12292_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_180_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14030_ _14030_/A vssd1 vssd1 vccd1 vccd1 _14030_/X sky130_fd_sc_hd__buf_8
X_11242_ _11892_/B _11242_/B vssd1 vssd1 vccd1 vccd1 _11245_/B sky130_fd_sc_hd__nand2_1
XFILLER_84_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11173_ _17805_/Q _11212_/B vssd1 vssd1 vccd1 vccd1 _11174_/C sky130_fd_sc_hd__or2_1
XFILLER_164_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10124_ _10124_/A _10124_/B vssd1 vssd1 vccd1 vccd1 _10124_/Y sky130_fd_sc_hd__nor2_1
XFILLER_164_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15981_ _18572_/Q _15980_/B _15980_/Y _15972_/X vssd1 vssd1 vccd1 vccd1 _18572_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_5620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17720_ _17720_/A vssd1 vssd1 vccd1 vccd1 _19004_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_76_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14932_ _14932_/A _14935_/B vssd1 vssd1 vccd1 vccd1 _14932_/Y sky130_fd_sc_hd__nand2_1
X_10055_ _09160_/B _10040_/A _09999_/A _09193_/C vssd1 vssd1 vccd1 vccd1 _10055_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17651_ _14597_/A _17649_/Y _17631_/X _17650_/Y _18975_/Q vssd1 vssd1 vccd1 vccd1
+ _17652_/B sky130_fd_sc_hd__a32o_1
XTAP_4963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14863_ _15156_/A _14989_/C vssd1 vssd1 vccd1 vccd1 _14875_/B sky130_fd_sc_hd__nor2_1
XTAP_4974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16602_ _16745_/A _16602_/B vssd1 vssd1 vccd1 vccd1 _16611_/B sky130_fd_sc_hd__nor2_1
XFILLER_17_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13814_ _18930_/Q _13772_/X _13654_/A _18927_/Q _13813_/X vssd1 vssd1 vccd1 vccd1
+ _13814_/X sky130_fd_sc_hd__a221o_1
XFILLER_21_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17582_ _17631_/A vssd1 vssd1 vccd1 vccd1 _17582_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_14794_ _14802_/B _14792_/X _14793_/X _14778_/X vssd1 vssd1 vccd1 vccd1 _18288_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_63_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_223_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_169_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16533_ _16538_/B _16531_/X _16532_/X _16519_/X vssd1 vssd1 vccd1 vccd1 _18702_/D
+ sky130_fd_sc_hd__o211a_1
X_13745_ _18333_/Q _13738_/X _13740_/X _13744_/X vssd1 vssd1 vccd1 vccd1 _13745_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_50_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_5_15_0_wb_clk_i clkbuf_4_7_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18102_/CLK
+ sky130_fd_sc_hd__clkbuf_2
X_10957_ _09408_/C _09709_/A _10956_/X _09987_/X vssd1 vssd1 vccd1 vccd1 _10957_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_17_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_182_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16464_ _16510_/A _16464_/B vssd1 vssd1 vccd1 vccd1 _16464_/Y sky130_fd_sc_hd__nand2_1
XFILLER_177_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13676_ _18549_/Q _13657_/X _13664_/X _18525_/Q vssd1 vssd1 vccd1 vccd1 _13676_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_182_1278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10888_ _10868_/X _10887_/X _10679_/X vssd1 vssd1 vccd1 vccd1 _10888_/X sky130_fd_sc_hd__o21a_1
X_18203_ _18203_/CLK _18203_/D vssd1 vssd1 vccd1 vccd1 _18203_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_223_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15415_ _15415_/A vssd1 vssd1 vccd1 vccd1 _15435_/S sky130_fd_sc_hd__clkbuf_2
X_19183_ _19183_/A _08999_/Y vssd1 vssd1 vccd1 vccd1 io_out[21] sky130_fd_sc_hd__ebufn_8
XFILLER_19_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12627_ _12627_/A _12627_/B vssd1 vssd1 vccd1 vccd1 _12628_/B sky130_fd_sc_hd__or2_1
X_16395_ _16689_/A _16452_/B vssd1 vssd1 vccd1 vccd1 _16407_/B sky130_fd_sc_hd__nor2_2
X_18134_ _18244_/CLK _18134_/D vssd1 vssd1 vccd1 vccd1 _18134_/Q sky130_fd_sc_hd__dfxtp_1
X_15346_ _15358_/A _15946_/B _15358_/C vssd1 vssd1 vccd1 vccd1 _15346_/X sky130_fd_sc_hd__or3_1
XFILLER_156_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12558_ _12557_/A _12557_/B _12529_/X vssd1 vssd1 vccd1 vccd1 _12558_/X sky130_fd_sc_hd__o21a_1
XFILLER_129_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18065_ _18072_/CLK _18065_/D vssd1 vssd1 vccd1 vccd1 _18065_/Q sky130_fd_sc_hd__dfxtp_1
X_11509_ _17872_/Q vssd1 vssd1 vccd1 vccd1 _11522_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_89_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15277_ _15277_/A _15277_/B vssd1 vssd1 vccd1 vccd1 _15286_/B sky130_fd_sc_hd__nor2_2
XFILLER_171_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12489_ _12492_/A _12487_/Y _12484_/X _12485_/Y vssd1 vssd1 vccd1 vccd1 _12490_/C
+ sky130_fd_sc_hd__o211ai_1
X_17016_ _17023_/B _17014_/X _17015_/X _16999_/X vssd1 vssd1 vccd1 vccd1 _18816_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_132_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14228_ _14332_/S _18994_/Q _14330_/B vssd1 vssd1 vccd1 vccd1 _14283_/A sky130_fd_sc_hd__or3_2
XFILLER_67_1333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14159_ _18770_/Q _14015_/X _14027_/X _18761_/Q _14158_/X vssd1 vssd1 vccd1 vccd1
+ _14159_/X sky130_fd_sc_hd__a221o_4
XFILLER_154_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_1208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18967_ _18967_/CLK _18967_/D vssd1 vssd1 vccd1 vccd1 _18967_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_47_wb_clk_i clkbuf_5_5_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18849_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17918_ _17919_/CLK _17918_/D vssd1 vssd1 vccd1 vccd1 _17918_/Q sky130_fd_sc_hd__dfxtp_1
X_18898_ _18899_/CLK _18898_/D vssd1 vssd1 vccd1 vccd1 _18898_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_152_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17849_ _19021_/CLK _17849_/D vssd1 vssd1 vccd1 vccd1 _17849_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_227_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_214_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_226_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_1304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_228_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_210_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09203_ _09203_/A _09203_/B _09203_/C _09203_/D vssd1 vssd1 vccd1 vccd1 _09204_/C
+ sky130_fd_sc_hd__and4_1
XFILLER_33_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_202_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09134_ _18809_/Q _18808_/Q _18807_/Q vssd1 vssd1 vccd1 vccd1 _09136_/C sky130_fd_sc_hd__or3_2
XFILLER_33_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09065_ _09072_/A _09069_/B _17826_/Q vssd1 vssd1 vccd1 vccd1 _09066_/A sky130_fd_sc_hd__and3_1
XFILLER_194_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_198_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09967_ _10388_/A vssd1 vssd1 vccd1 vccd1 _14260_/B sky130_fd_sc_hd__buf_4
XTAP_4204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_218_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09898_ _09924_/A vssd1 vssd1 vccd1 vccd1 _10600_/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_217_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11860_ _11860_/A _11860_/B vssd1 vssd1 vccd1 vccd1 _11860_/Y sky130_fd_sc_hd__nor2_1
XTAP_2824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10811_ _10811_/A _10811_/B vssd1 vssd1 vccd1 vccd1 _10811_/X sky130_fd_sc_hd__or2_1
XFILLER_32_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11791_ _11753_/A _11654_/B _11404_/B _11593_/A _11737_/B vssd1 vssd1 vccd1 vccd1
+ _11791_/X sky130_fd_sc_hd__o2111a_1
XTAP_2868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13530_ _13731_/A vssd1 vssd1 vccd1 vccd1 _13531_/A sky130_fd_sc_hd__buf_6
X_10742_ _09103_/C _09098_/D _10763_/S vssd1 vssd1 vccd1 vccd1 _10743_/B sky130_fd_sc_hd__mux2_1
XFILLER_201_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13461_ _13467_/A _13461_/B vssd1 vssd1 vccd1 vccd1 _18154_/D sky130_fd_sc_hd__nor2_1
X_10673_ _10864_/A _10679_/A _10649_/X _10672_/X vssd1 vssd1 vccd1 vccd1 _10673_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_41_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15200_ _15206_/B _15198_/X _15199_/X _15187_/X vssd1 vssd1 vccd1 vccd1 _18387_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_139_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12412_ _12412_/A _12412_/B vssd1 vssd1 vccd1 vccd1 _12414_/C sky130_fd_sc_hd__nor2_1
X_16180_ _16935_/A vssd1 vssd1 vccd1 vccd1 _16773_/B sky130_fd_sc_hd__buf_4
XFILLER_138_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13392_ _18121_/Q _11040_/X _11035_/B _13381_/X _13383_/A vssd1 vssd1 vccd1 vccd1
+ _18121_/D sky130_fd_sc_hd__o2111a_1
X_15131_ _15252_/A vssd1 vssd1 vccd1 vccd1 _15182_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_166_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12343_ _11478_/A _11478_/B _12342_/X _12318_/X vssd1 vssd1 vccd1 vccd1 _17887_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_177_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15062_ _15061_/B _15060_/X _15061_/Y _15046_/X vssd1 vssd1 vccd1 vccd1 _18353_/D
+ sky130_fd_sc_hd__o211a_1
X_12274_ _12274_/A _12276_/C vssd1 vssd1 vccd1 vccd1 _12274_/Y sky130_fd_sc_hd__nor2_1
XFILLER_177_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_141_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11225_ _11237_/C vssd1 vssd1 vccd1 vccd1 _11232_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_49_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14013_ _14013_/A vssd1 vssd1 vccd1 vccd1 _18167_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_153_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18821_ _18821_/CLK _18821_/D vssd1 vssd1 vccd1 vccd1 _18821_/Q sky130_fd_sc_hd__dfxtp_4
X_11156_ _11156_/A vssd1 vssd1 vccd1 vccd1 _17803_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_67_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_191_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10107_ _12068_/A _10940_/A _10094_/X _10100_/X _10106_/X vssd1 vssd1 vccd1 vccd1
+ _10107_/X sky130_fd_sc_hd__a311o_1
X_18752_ _18752_/CLK _18752_/D vssd1 vssd1 vccd1 vccd1 _18752_/Q sky130_fd_sc_hd__dfxtp_2
X_15964_ _15984_/A _15964_/B _15964_/C vssd1 vssd1 vccd1 vccd1 _15964_/X sky130_fd_sc_hd__or3_1
XTAP_5450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11087_ _11313_/B _11001_/C _11091_/S vssd1 vssd1 vccd1 vccd1 _11088_/A sky130_fd_sc_hd__mux2_1
XFILLER_209_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17703_ _17703_/A vssd1 vssd1 vccd1 vccd1 _18988_/D sky130_fd_sc_hd__clkbuf_1
XTAP_5483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10038_ _10007_/B _10038_/B vssd1 vssd1 vccd1 vccd1 _10039_/A sky130_fd_sc_hd__and2b_1
X_14915_ _14915_/A vssd1 vssd1 vccd1 vccd1 _16431_/A sky130_fd_sc_hd__buf_12
X_18683_ _18683_/CLK _18683_/D vssd1 vssd1 vccd1 vccd1 _18683_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_5494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15895_ _15900_/B _15893_/X _15894_/X _15881_/X vssd1 vssd1 vccd1 vccd1 _18552_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_4760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_209_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17634_ _17634_/A vssd1 vssd1 vccd1 vccd1 _18971_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_184_1307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14846_ _14872_/A _14849_/B vssd1 vssd1 vccd1 vccd1 _14846_/Y sky130_fd_sc_hd__nand2_1
XFILLER_1_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_208_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_184_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_223_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17565_ _17565_/A vssd1 vssd1 vccd1 vccd1 _18954_/D sky130_fd_sc_hd__clkbuf_1
X_14777_ _14814_/A _14777_/B vssd1 vssd1 vccd1 vccd1 _14777_/Y sky130_fd_sc_hd__nand2_1
X_11989_ _12027_/C _13434_/C vssd1 vssd1 vccd1 vccd1 _11990_/C sky130_fd_sc_hd__nor2_1
X_16516_ _16578_/A vssd1 vssd1 vccd1 vccd1 _16650_/B sky130_fd_sc_hd__clkbuf_2
X_13728_ _18237_/Q _13544_/A _13718_/X _13727_/X vssd1 vssd1 vccd1 vccd1 _13728_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_225_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_204_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17496_ _17509_/A _17501_/B vssd1 vssd1 vccd1 vccd1 _17496_/Y sky130_fd_sc_hd__nand2_1
XFILLER_220_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_165_wb_clk_i clkbuf_5_10_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18072_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_108_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_231_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19235_ _19235_/A _08945_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[35] sky130_fd_sc_hd__ebufn_8
X_16447_ _16447_/A _16450_/B vssd1 vssd1 vccd1 vccd1 _16447_/Y sky130_fd_sc_hd__nand2_1
X_13659_ _18969_/Q _13705_/A _13706_/A _18951_/Q vssd1 vssd1 vccd1 vccd1 _13659_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_176_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19166_ _19166_/A _09030_/Y vssd1 vssd1 vccd1 vccd1 io_out[4] sky130_fd_sc_hd__ebufn_8
XFILLER_121_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16378_ _16392_/A _16378_/B vssd1 vssd1 vccd1 vccd1 _16378_/Y sky130_fd_sc_hd__nand2_1
XFILLER_9_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18117_ _18126_/CLK _18117_/D vssd1 vssd1 vccd1 vccd1 _18117_/Q sky130_fd_sc_hd__dfxtp_1
X_15329_ _15931_/A _15393_/B vssd1 vssd1 vccd1 vccd1 _15339_/B sky130_fd_sc_hd__nor2_2
XFILLER_8_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_219_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18048_ _18052_/CLK _18048_/D vssd1 vssd1 vccd1 vccd1 _18048_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_99_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09821_ _18113_/Q vssd1 vssd1 vccd1 vccd1 _09844_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_87_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09752_ _09752_/A _09752_/B vssd1 vssd1 vccd1 vccd1 _09753_/B sky130_fd_sc_hd__or2_1
XFILLER_80_1352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_230_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09683_ _10085_/S vssd1 vssd1 vccd1 vccd1 _09683_/X sky130_fd_sc_hd__buf_6
XFILLER_41_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_215_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_215_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_223_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_210_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_183_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_183_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09117_ _18758_/Q _18757_/Q _18756_/Q vssd1 vssd1 vccd1 vccd1 _09119_/C sky130_fd_sc_hd__or3_4
XFILLER_135_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09048_ _09052_/A vssd1 vssd1 vccd1 vccd1 _09048_/Y sky130_fd_sc_hd__inv_2
XFILLER_164_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11010_ _11181_/A _17806_/Q _17808_/Q vssd1 vssd1 vccd1 vccd1 _11011_/D sky130_fd_sc_hd__nand3b_1
XFILLER_104_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_219_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_219_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_40 _10089_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12961_ _12961_/A _12961_/B vssd1 vssd1 vccd1 vccd1 _12969_/B sky130_fd_sc_hd__and2_1
XFILLER_79_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_51 _10648_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_218_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14700_ _14753_/A _14700_/B vssd1 vssd1 vccd1 vccd1 _14700_/Y sky130_fd_sc_hd__nand2_1
XINSDIODE2_62 _17747_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_73 _13576_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11912_ _17977_/Q vssd1 vssd1 vccd1 vccd1 _12982_/A sky130_fd_sc_hd__buf_6
X_15680_ _15691_/A _15683_/B vssd1 vssd1 vccd1 vccd1 _15680_/Y sky130_fd_sc_hd__nand2_1
XINSDIODE2_84 _13619_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XINSDIODE2_95 _13721_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12892_ _12895_/C _12892_/B vssd1 vssd1 vccd1 vccd1 _17960_/D sky130_fd_sc_hd__nor2_1
XTAP_2621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14631_ _17541_/A vssd1 vssd1 vccd1 vccd1 _14681_/A sky130_fd_sc_hd__buf_2
XTAP_3388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11843_ _11848_/A _11843_/B vssd1 vssd1 vccd1 vccd1 _11844_/B sky130_fd_sc_hd__nor2_1
XFILLER_54_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17350_ _17349_/B _17347_/X _17349_/Y _17341_/X vssd1 vssd1 vccd1 vccd1 _18899_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_2687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14562_ _18236_/Q _14559_/B _14559_/Y _14561_/X vssd1 vssd1 vccd1 vccd1 _18236_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_13_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11774_ _11758_/X _11766_/X _11773_/X vssd1 vssd1 vccd1 vccd1 _11774_/Y sky130_fd_sc_hd__o21ai_1
XTAP_1964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16301_ _18682_/Q _18646_/Q _16304_/S vssd1 vssd1 vccd1 vccd1 _16301_/X sky130_fd_sc_hd__mux2_1
XFILLER_202_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_213_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13513_ _13513_/A vssd1 vssd1 vccd1 vccd1 _13582_/A sky130_fd_sc_hd__buf_6
XFILLER_201_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10725_ _10753_/A _10718_/X _10724_/X _10616_/Y vssd1 vssd1 vccd1 vccd1 _10725_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_1997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17281_ _18918_/Q _18882_/Q _17298_/S vssd1 vssd1 vccd1 vccd1 _17281_/X sky130_fd_sc_hd__mux2_1
XFILLER_144_1368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14493_ _17420_/A vssd1 vssd1 vccd1 vccd1 _14502_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_13_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19020_ _19026_/CLK _19020_/D vssd1 vssd1 vccd1 vccd1 _19020_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_41_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16232_ _16672_/A _16358_/C vssd1 vssd1 vccd1 vccd1 _16243_/B sky130_fd_sc_hd__nor2_1
X_13444_ _13444_/A _11364_/B vssd1 vssd1 vccd1 vccd1 _13444_/X sky130_fd_sc_hd__or2b_1
XFILLER_186_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10656_ _18122_/Q _10656_/B vssd1 vssd1 vccd1 vccd1 _10721_/A sky130_fd_sc_hd__xnor2_4
XFILLER_16_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16163_ _16160_/B _16159_/X _16160_/Y _16162_/X vssd1 vssd1 vccd1 vccd1 _18614_/D
+ sky130_fd_sc_hd__o211a_1
X_10587_ _09294_/C _09299_/B _09304_/D _09299_/D _10096_/S _09682_/A vssd1 vssd1 vccd1
+ vccd1 _10587_/X sky130_fd_sc_hd__mux4_1
X_13375_ _13375_/A _13375_/B _13375_/C _13394_/D vssd1 vssd1 vccd1 vccd1 _13379_/B
+ sky130_fd_sc_hd__nor4b_4
XFILLER_155_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15114_ _18403_/Q _18367_/Q _15121_/S vssd1 vssd1 vccd1 vccd1 _15114_/X sky130_fd_sc_hd__mux2_1
X_12326_ _12329_/B _12327_/A _12327_/B _12329_/A vssd1 vssd1 vccd1 vccd1 _12330_/A
+ sky130_fd_sc_hd__a31o_1
X_16094_ _16173_/A vssd1 vssd1 vccd1 vccd1 _16113_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_181_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_177_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15045_ _15058_/A _15049_/B vssd1 vssd1 vccd1 vccd1 _15045_/Y sky130_fd_sc_hd__nand2_1
X_12257_ _12257_/A vssd1 vssd1 vccd1 vccd1 _13066_/B sky130_fd_sc_hd__buf_8
XFILLER_141_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11208_ _11209_/A _11209_/B vssd1 vssd1 vccd1 vccd1 _11210_/B sky130_fd_sc_hd__nand2_1
X_12188_ _12444_/B vssd1 vssd1 vccd1 vccd1 _12470_/B sky130_fd_sc_hd__buf_2
XFILLER_64_1347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_218_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_214_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18804_ _18806_/CLK _18804_/D vssd1 vssd1 vccd1 vccd1 _18804_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_95_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11139_ _17801_/Q vssd1 vssd1 vccd1 vccd1 _11498_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_96_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_231_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16996_ _16998_/B _16994_/X _16995_/Y _16964_/X vssd1 vssd1 vccd1 vccd1 _18811_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_110_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15947_ _16273_/A vssd1 vssd1 vccd1 vccd1 _16028_/A sky130_fd_sc_hd__clkbuf_2
X_18735_ _18738_/CLK _18735_/D vssd1 vssd1 vccd1 vccd1 _18735_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_114_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18666_ _18683_/CLK _18666_/D vssd1 vssd1 vccd1 vccd1 _18666_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_224_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15878_ _16030_/A _15892_/B vssd1 vssd1 vccd1 vccd1 _15890_/B sky130_fd_sc_hd__nor2_2
XTAP_4590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14829_ _15266_/A _14841_/B vssd1 vssd1 vccd1 vccd1 _14838_/B sky130_fd_sc_hd__nor2_2
XFILLER_63_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17617_ _17616_/Y _17552_/X _18966_/Q vssd1 vssd1 vccd1 vccd1 _17617_/X sky130_fd_sc_hd__a21o_1
XFILLER_97_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18597_ _18608_/CLK _18597_/D vssd1 vssd1 vccd1 vccd1 _18597_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_36_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_225_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_229_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17548_ _17602_/A _17687_/A vssd1 vssd1 vccd1 vccd1 _17548_/Y sky130_fd_sc_hd__nor2_1
XFILLER_225_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_1318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17479_ _18932_/Q _17477_/B _17477_/Y _17478_/X vssd1 vssd1 vccd1 vccd1 _18932_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_221_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_225_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19218_ _19218_/A _08962_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[18] sky130_fd_sc_hd__ebufn_8
XFILLER_20_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_220_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19149_ _19149_/A _09038_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[19] sky130_fd_sc_hd__ebufn_8
XFILLER_117_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_5_8_0_wb_clk_i clkbuf_5_9_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_5_8_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_160_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_62_wb_clk_i clkbuf_5_20_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18701_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_120_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09804_ _09743_/A _10675_/A _09803_/X vssd1 vssd1 vccd1 vccd1 _09805_/B sky130_fd_sc_hd__o21a_1
XFILLER_86_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09735_ _19027_/Q _10618_/A vssd1 vssd1 vccd1 vccd1 _09735_/Y sky130_fd_sc_hd__nand2_1
XFILLER_101_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_189_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_216_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_227_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09666_ _09664_/A _09630_/B _09665_/X vssd1 vssd1 vccd1 vccd1 _09667_/B sky130_fd_sc_hd__o21a_1
XFILLER_27_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_216_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_199_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09597_ _09588_/X _09726_/A _09596_/X vssd1 vssd1 vccd1 vccd1 _09611_/A sky130_fd_sc_hd__a21o_1
XTAP_1227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_230_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_208_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_204_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10510_ _10443_/A _10508_/X _10509_/X _10183_/A _10454_/X vssd1 vssd1 vccd1 vccd1
+ _10510_/X sky130_fd_sc_hd__a221o_2
X_11490_ _12336_/B vssd1 vssd1 vccd1 vccd1 _11490_/Y sky130_fd_sc_hd__inv_2
XFILLER_7_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10441_ _10441_/A _10441_/B vssd1 vssd1 vccd1 vccd1 _12031_/A sky130_fd_sc_hd__or2_4
XFILLER_148_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13160_ _13164_/A _18039_/Q vssd1 vssd1 vccd1 vccd1 _13161_/A sky130_fd_sc_hd__and2_1
X_10372_ _10605_/C _10365_/X _10366_/X _10371_/X vssd1 vssd1 vccd1 vccd1 _10372_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_200_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12111_ _12112_/B _12112_/C _12112_/A vssd1 vssd1 vccd1 vccd1 _12111_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_123_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13091_ _13091_/A vssd1 vssd1 vccd1 vccd1 _18007_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_151_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12042_ _12042_/A _12042_/B vssd1 vssd1 vccd1 vccd1 _12043_/B sky130_fd_sc_hd__nor2_1
XFILLER_123_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_215_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16850_ _16850_/A vssd1 vssd1 vccd1 vccd1 _17446_/A sky130_fd_sc_hd__buf_4
XFILLER_215_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15801_ _18565_/Q _18529_/Q _15809_/S vssd1 vssd1 vccd1 vccd1 _15801_/X sky130_fd_sc_hd__mux2_1
XFILLER_1_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_219_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16781_ _16871_/A vssd1 vssd1 vccd1 vccd1 _16781_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_1_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13993_ _18577_/Q _13760_/A _13781_/A _18568_/Q vssd1 vssd1 vccd1 vccd1 _13993_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_65_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_219_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_218_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18520_ _18546_/CLK _18520_/D vssd1 vssd1 vccd1 vccd1 _18520_/Q sky130_fd_sc_hd__dfxtp_2
X_15732_ _16030_/A _15745_/B vssd1 vssd1 vccd1 vccd1 _15743_/B sky130_fd_sc_hd__nor2_2
XFILLER_65_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12944_ _13049_/A _12944_/B vssd1 vssd1 vccd1 vccd1 _12945_/A sky130_fd_sc_hd__and2_1
XFILLER_74_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18451_ _18467_/CLK _18451_/D vssd1 vssd1 vccd1 vccd1 _18451_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_206_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15663_ _15661_/B _15660_/X _15661_/Y _15662_/X vssd1 vssd1 vccd1 vccd1 _18494_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_45_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_222_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_209_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12875_ _12824_/A _12877_/C _12874_/X vssd1 vssd1 vccd1 vccd1 _12875_/Y sky130_fd_sc_hd__o21ai_1
XTAP_3185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17402_ _18949_/Q _18913_/Q _17406_/S vssd1 vssd1 vccd1 vccd1 _17402_/X sky130_fd_sc_hd__mux2_1
X_14614_ _14354_/X _14608_/X _14612_/X _14613_/Y _11822_/X vssd1 vssd1 vccd1 vccd1
+ _18246_/D sky130_fd_sc_hd__o311a_1
XTAP_2473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18382_ _18406_/CLK _18382_/D vssd1 vssd1 vccd1 vccd1 _18382_/Q sky130_fd_sc_hd__dfxtp_2
X_11826_ _11826_/A _11826_/B _11826_/C vssd1 vssd1 vccd1 vccd1 _11826_/X sky130_fd_sc_hd__or3_1
XTAP_2484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15594_ _15633_/A _15594_/B vssd1 vssd1 vccd1 vccd1 _15594_/Y sky130_fd_sc_hd__nand2_1
XTAP_1750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_202_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_109_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_159_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17333_ _18894_/Q _17336_/B _17332_/X _17324_/X vssd1 vssd1 vccd1 vccd1 _18894_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_159_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14545_ _14606_/A _14545_/B vssd1 vssd1 vccd1 vccd1 _14545_/Y sky130_fd_sc_hd__nand2_1
XTAP_1783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11757_ _11757_/A _11797_/A vssd1 vssd1 vccd1 vccd1 _11757_/Y sky130_fd_sc_hd__nand2_1
XTAP_1794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_222_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17264_ _17263_/B _17262_/X _17263_/Y _17260_/X vssd1 vssd1 vccd1 vccd1 _18878_/D
+ sky130_fd_sc_hd__o211a_1
X_10708_ _12094_/A _10700_/X _10704_/X _10707_/Y vssd1 vssd1 vccd1 vccd1 _10708_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_147_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14476_ _18213_/Q _14480_/B vssd1 vssd1 vccd1 vccd1 _14477_/A sky130_fd_sc_hd__and2_1
X_11688_ _11703_/A _17850_/Q vssd1 vssd1 vccd1 vccd1 _11700_/A sky130_fd_sc_hd__nor2_1
X_19003_ _19004_/CLK _19003_/D vssd1 vssd1 vccd1 vccd1 _19003_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16215_ _18662_/Q _18626_/Q _16215_/S vssd1 vssd1 vccd1 vccd1 _16215_/X sky130_fd_sc_hd__mux2_1
X_13427_ _13427_/A vssd1 vssd1 vccd1 vccd1 _13447_/B sky130_fd_sc_hd__inv_2
X_17195_ _18898_/Q _18862_/Q _17199_/S vssd1 vssd1 vccd1 vccd1 _17195_/X sky130_fd_sc_hd__mux2_1
X_10639_ _10766_/A vssd1 vssd1 vccd1 vccd1 _10679_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_31_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16146_ _16216_/A vssd1 vssd1 vccd1 vccd1 _16202_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_161_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13358_ _14422_/A _14383_/C _14507_/B vssd1 vssd1 vccd1 vccd1 _14384_/B sky130_fd_sc_hd__a21oi_2
XFILLER_6_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12309_ _12327_/A _12327_/B vssd1 vssd1 vccd1 vccd1 _12333_/C sky130_fd_sc_hd__nand2_1
X_16077_ _16212_/A vssd1 vssd1 vccd1 vccd1 _16130_/A sky130_fd_sc_hd__clkbuf_2
X_13289_ _18017_/Q _18016_/Q _18019_/Q _18018_/Q vssd1 vssd1 vccd1 vccd1 _13291_/C
+ sky130_fd_sc_hd__or4_1
XFILLER_5_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15028_ _15064_/A vssd1 vssd1 vccd1 vccd1 _15085_/B sky130_fd_sc_hd__buf_2
XFILLER_102_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_229_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_229_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16979_ _16975_/A _16978_/X _18807_/Q vssd1 vssd1 vccd1 vccd1 _16979_/Y sky130_fd_sc_hd__o21bai_1
XFILLER_7_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput3 io_in[25] vssd1 vssd1 vccd1 vccd1 input3/X sky130_fd_sc_hd__clkbuf_1
XFILLER_49_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09520_ _19000_/Q vssd1 vssd1 vccd1 vccd1 _14319_/S sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_83_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18718_ _18719_/CLK _18718_/D vssd1 vssd1 vccd1 vccd1 _18718_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_225_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_180_wb_clk_i clkbuf_5_10_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _19004_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_149_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_224_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09451_ _09339_/A _09443_/Y _09420_/X _09450_/Y vssd1 vssd1 vccd1 vccd1 _09451_/X
+ sky130_fd_sc_hd__a22o_2
XFILLER_24_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18649_ _18650_/CLK _18649_/D vssd1 vssd1 vccd1 vccd1 _18649_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_224_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09382_ _18389_/Q _18388_/Q _18387_/Q vssd1 vssd1 vccd1 vccd1 _09386_/A sky130_fd_sc_hd__or3_4
XFILLER_149_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_123_1216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_137_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_119_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_195_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_69_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_117_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_1266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09718_ _09712_/X _09713_/X _09714_/X _09715_/X _10944_/S _09689_/X vssd1 vssd1 vccd1
+ vccd1 _09718_/X sky130_fd_sc_hd__mux4_1
XFILLER_28_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10990_ _10990_/A vssd1 vssd1 vccd1 vccd1 _10990_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_56_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09649_ _09649_/A _09649_/B _09704_/A vssd1 vssd1 vccd1 vccd1 _09649_/X sky130_fd_sc_hd__or3_2
XFILLER_216_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_203_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_231_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_215_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12660_ _17934_/Q vssd1 vssd1 vccd1 vccd1 _12662_/A sky130_fd_sc_hd__clkinv_2
XFILLER_169_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11611_ _17856_/Q _11624_/B vssd1 vssd1 vccd1 vccd1 _11623_/B sky130_fd_sc_hd__nor2_1
XFILLER_208_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12591_ _12591_/A vssd1 vssd1 vccd1 vccd1 _12591_/X sky130_fd_sc_hd__buf_2
XFILLER_212_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_204_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14330_ _14330_/A _14330_/B vssd1 vssd1 vccd1 vccd1 _14330_/Y sky130_fd_sc_hd__nor2_1
XFILLER_184_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11542_ _11921_/B _11542_/B vssd1 vssd1 vccd1 vccd1 _13518_/A sky130_fd_sc_hd__and2_2
XFILLER_195_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_1338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14261_ _14260_/A _14259_/Y _14260_/Y _14272_/A vssd1 vssd1 vccd1 vccd1 _14261_/X
+ sky130_fd_sc_hd__o211a_1
X_11473_ _17888_/Q vssd1 vssd1 vccd1 vccd1 _11473_/Y sky130_fd_sc_hd__inv_2
XFILLER_7_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16000_ _16000_/A _16003_/B vssd1 vssd1 vccd1 vccd1 _16000_/Y sky130_fd_sc_hd__nand2_1
XFILLER_171_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13212_ _17661_/A vssd1 vssd1 vccd1 vccd1 _13257_/A sky130_fd_sc_hd__buf_2
XFILLER_137_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10424_ _12039_/A _10415_/Y _10419_/Y _10421_/Y _10533_/B vssd1 vssd1 vccd1 vccd1
+ _10424_/X sky130_fd_sc_hd__a311o_1
XFILLER_139_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14192_ _18208_/Q _14233_/A _18209_/Q vssd1 vssd1 vccd1 vccd1 _14192_/X sky130_fd_sc_hd__a21o_1
XFILLER_87_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13143_ _13151_/A _18031_/Q vssd1 vssd1 vccd1 vccd1 _13144_/A sky130_fd_sc_hd__and2_1
X_10355_ _09153_/A _09143_/B _09148_/C _10722_/A _09958_/A _09948_/A vssd1 vssd1 vccd1
+ vccd1 _10356_/B sky130_fd_sc_hd__mux4_1
XFILLER_87_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_215_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10286_ _09203_/C _09193_/C _10286_/S vssd1 vssd1 vccd1 vccd1 _10286_/X sky130_fd_sc_hd__mux2_1
XTAP_819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13074_ _14533_/A vssd1 vssd1 vccd1 vccd1 _13074_/X sky130_fd_sc_hd__clkbuf_2
X_17951_ _17954_/CLK _17951_/D vssd1 vssd1 vccd1 vccd1 _17951_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_105_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_215_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16902_ _17168_/A vssd1 vssd1 vccd1 vccd1 _16957_/A sky130_fd_sc_hd__buf_2
X_12025_ _12025_/A _12025_/B _12026_/B _12025_/D vssd1 vssd1 vccd1 vccd1 _12027_/B
+ sky130_fd_sc_hd__and4_4
X_17882_ _17883_/CLK _17882_/D vssd1 vssd1 vccd1 vccd1 _17882_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_104_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_215_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16833_ _16884_/A _16833_/B vssd1 vssd1 vccd1 vccd1 _16833_/Y sky130_fd_sc_hd__nand2_1
XFILLER_66_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16764_ _16813_/A _16769_/B vssd1 vssd1 vccd1 vccd1 _16764_/Y sky130_fd_sc_hd__nand2_1
X_13976_ _18274_/Q _13733_/X _13972_/X _13975_/X vssd1 vssd1 vccd1 vccd1 _13976_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_65_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_219_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18503_ _18504_/CLK _18503_/D vssd1 vssd1 vccd1 vccd1 _18503_/Q sky130_fd_sc_hd__dfxtp_4
X_15715_ _15751_/A _15719_/B vssd1 vssd1 vccd1 vccd1 _15715_/Y sky130_fd_sc_hd__nand2_1
XFILLER_18_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_207_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12927_ _12927_/A _12931_/A vssd1 vssd1 vccd1 vccd1 _12927_/Y sky130_fd_sc_hd__nand2_1
X_16695_ _16695_/A _16699_/B vssd1 vssd1 vccd1 vccd1 _16695_/Y sky130_fd_sc_hd__nand2_1
XFILLER_146_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15646_ _15651_/B _15642_/X _15645_/Y _15640_/X vssd1 vssd1 vccd1 vccd1 _18490_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_222_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18434_ _18434_/CLK _18434_/D vssd1 vssd1 vccd1 vccd1 _18434_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_179_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12858_ _17948_/Q _12816_/X _12851_/B _17950_/Q vssd1 vssd1 vccd1 vccd1 _12859_/B
+ sky130_fd_sc_hd__a31o_1
XTAP_2270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18365_ _18392_/CLK _18365_/D vssd1 vssd1 vccd1 vccd1 _18365_/Q sky130_fd_sc_hd__dfxtp_2
X_11809_ _11781_/A _11780_/Y _11800_/X _11869_/B vssd1 vssd1 vccd1 vccd1 _11809_/X
+ sky130_fd_sc_hd__a211o_1
X_15577_ _18511_/Q _18475_/Q _15586_/S vssd1 vssd1 vccd1 vccd1 _15577_/X sky130_fd_sc_hd__mux2_1
XTAP_1580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12789_ _13085_/A _12788_/Y _12786_/B vssd1 vssd1 vccd1 vccd1 _12789_/X sky130_fd_sc_hd__o21a_1
XFILLER_221_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17316_ _17458_/A _17351_/B vssd1 vssd1 vccd1 vccd1 _17327_/B sky130_fd_sc_hd__nor2_1
XFILLER_187_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14528_ _17415_/B _14690_/B vssd1 vssd1 vccd1 vccd1 _14545_/B sky130_fd_sc_hd__nor2_2
XFILLER_30_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18296_ _18296_/CLK _18296_/D vssd1 vssd1 vccd1 vccd1 _18296_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_202_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17247_ _17247_/A vssd1 vssd1 vccd1 vccd1 _17262_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_31_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19128__99 vssd1 vssd1 vccd1 vccd1 _19128__99/HI _19236_/A sky130_fd_sc_hd__conb_1
X_14459_ _14279_/A _17709_/B _12764_/X vssd1 vssd1 vccd1 vccd1 _14459_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_134_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17178_ _17180_/B _17176_/X _17177_/Y _17161_/X vssd1 vssd1 vccd1 vccd1 _18856_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_155_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16129_ _18606_/Q _16132_/B _16128_/X _16120_/X vssd1 vssd1 vccd1 vccd1 _18606_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_6_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_1334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08951_ _08954_/A vssd1 vssd1 vccd1 vccd1 _08951_/Y sky130_fd_sc_hd__inv_2
XFILLER_103_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_229_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09503_ _18201_/Q _09503_/B vssd1 vssd1 vccd1 vccd1 _14445_/B sky130_fd_sc_hd__or2_1
XFILLER_77_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_225_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_213_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09434_ _09434_/A vssd1 vssd1 vccd1 vccd1 _18150_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_53_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_205_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09365_ _09365_/A _09365_/B _09365_/C _09365_/D vssd1 vssd1 vccd1 vccd1 _09371_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_212_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_221_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_205_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09296_ _18503_/Q _18502_/Q _18501_/Q vssd1 vssd1 vccd1 vccd1 _09299_/B sky130_fd_sc_hd__or3_4
XFILLER_165_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10140_ _10140_/A _10160_/B vssd1 vssd1 vccd1 vccd1 _10141_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10071_ _09237_/A _09227_/B _09232_/C _09237_/C _10060_/X _10025_/X vssd1 vssd1 vccd1
+ vccd1 _10071_/X sky130_fd_sc_hd__mux4_1
XTAP_5824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_1216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13830_ _11957_/B _13634_/X _13712_/X _13829_/X vssd1 vssd1 vccd1 vccd1 _13830_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_47_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13761_ _18504_/Q _13847_/A _13654_/A _18495_/Q vssd1 vssd1 vccd1 vccd1 _13761_/X
+ sky130_fd_sc_hd__a22o_1
XINSDIODE2_209 _13546_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10973_ _17941_/Q vssd1 vssd1 vccd1 vccd1 _13418_/B sky130_fd_sc_hd__inv_2
XFILLER_46_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15500_ _15511_/A _15500_/B vssd1 vssd1 vccd1 vccd1 _15500_/Y sky130_fd_sc_hd__nand2_1
XFILLER_71_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12712_ _17938_/Q _12707_/X _17939_/Q vssd1 vssd1 vccd1 vccd1 _12713_/B sky130_fd_sc_hd__o21ai_1
X_16480_ _18726_/Q _18690_/Q _16490_/S vssd1 vssd1 vccd1 vccd1 _16480_/X sky130_fd_sc_hd__mux2_1
XPHY_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_231_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13692_ _18597_/Q _13544_/A _13688_/X _13691_/X vssd1 vssd1 vccd1 vccd1 _13692_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_15_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_204_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15431_ _15445_/A _15431_/B vssd1 vssd1 vccd1 vccd1 _15431_/Y sky130_fd_sc_hd__nand2_1
XFILLER_43_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12643_ _17929_/Q vssd1 vssd1 vccd1 vccd1 _12646_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_43_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18150_ _18251_/CLK _18150_/D vssd1 vssd1 vccd1 vccd1 _18150_/Q sky130_fd_sc_hd__dfxtp_1
X_15362_ _15373_/A _15366_/B vssd1 vssd1 vccd1 vccd1 _15362_/Y sky130_fd_sc_hd__nand2_1
XFILLER_197_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_212_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12574_ _17924_/Q _12574_/B vssd1 vssd1 vccd1 vccd1 _12575_/B sky130_fd_sc_hd__nor2_1
XFILLER_106_1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17101_ _17152_/A _17105_/B vssd1 vssd1 vccd1 vccd1 _17101_/Y sky130_fd_sc_hd__nand2_1
XFILLER_178_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14313_ _13409_/X _14306_/X _14310_/Y _14312_/X vssd1 vssd1 vccd1 vccd1 _14313_/X
+ sky130_fd_sc_hd__o22a_1
X_18081_ _18087_/CLK _18081_/D vssd1 vssd1 vccd1 vccd1 _18081_/Q sky130_fd_sc_hd__dfxtp_1
X_11525_ _11828_/A _11525_/B vssd1 vssd1 vccd1 vccd1 _11701_/A sky130_fd_sc_hd__and2_1
X_15293_ _18182_/Q vssd1 vssd1 vccd1 vccd1 _16566_/A sky130_fd_sc_hd__buf_6
XFILLER_7_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17032_ _17032_/A _17035_/B vssd1 vssd1 vccd1 vccd1 _17032_/Y sky130_fd_sc_hd__nand2_1
XFILLER_116_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14244_ _14300_/A vssd1 vssd1 vccd1 vccd1 _14244_/X sky130_fd_sc_hd__clkbuf_2
X_11456_ _17887_/Q vssd1 vssd1 vccd1 vccd1 _11459_/A sky130_fd_sc_hd__inv_2
XFILLER_171_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10407_ _10314_/X _10336_/X _10360_/X _10405_/X _10406_/Y vssd1 vssd1 vccd1 vccd1
+ _13411_/A sky130_fd_sc_hd__o41a_1
X_14175_ _18683_/Q _13525_/X _14027_/A _18689_/Q vssd1 vssd1 vccd1 vccd1 _14175_/X
+ sky130_fd_sc_hd__a22o_1
X_11387_ _11323_/A _12299_/B _11339_/C vssd1 vssd1 vccd1 vccd1 _11388_/B sky130_fd_sc_hd__o21a_1
XFILLER_113_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13126_ _13126_/A vssd1 vssd1 vccd1 vccd1 _18022_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_152_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10338_ _10338_/A _10338_/B vssd1 vssd1 vccd1 vccd1 _10338_/X sky130_fd_sc_hd__and2_1
XFILLER_3_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18983_ _18986_/CLK _18983_/D vssd1 vssd1 vccd1 vccd1 _18983_/Q sky130_fd_sc_hd__dfxtp_2
Xclkbuf_leaf_119_wb_clk_i clkbuf_5_30_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18473_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_139_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13057_ _13375_/C _12776_/X _13056_/X _13037_/X vssd1 vssd1 vccd1 vccd1 _17996_/D
+ sky130_fd_sc_hd__o211a_1
X_17934_ _18902_/CLK _17934_/D vssd1 vssd1 vccd1 vccd1 _17934_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_112_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10269_ _11924_/A _10267_/X _10918_/S vssd1 vssd1 vccd1 vccd1 _10270_/C sky130_fd_sc_hd__a21o_1
XFILLER_6_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_1204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12008_ _12007_/A _12026_/C _12026_/D _12007_/Y vssd1 vssd1 vccd1 vccd1 _12009_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_121_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17865_ _19032_/CLK _17865_/D vssd1 vssd1 vccd1 vccd1 _17865_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_78_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_227_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16816_ _18773_/Q _16815_/B _16815_/Y _16800_/X vssd1 vssd1 vccd1 vccd1 _18773_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_213_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17796_ _17806_/CLK _17796_/D vssd1 vssd1 vccd1 vccd1 _17796_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_47_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_228_1302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13959_ _18646_/Q _13723_/X _13743_/X _18628_/Q vssd1 vssd1 vccd1 vccd1 _13959_/X
+ sky130_fd_sc_hd__a22o_1
X_16747_ _18792_/Q _18756_/Q _16762_/S vssd1 vssd1 vccd1 vccd1 _16747_/X sky130_fd_sc_hd__mux2_1
XFILLER_47_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_179_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16678_ _16678_/A _16678_/B _16716_/C vssd1 vssd1 vccd1 vccd1 _16678_/X sky130_fd_sc_hd__or3_1
XFILLER_222_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18417_ _18423_/CLK _18417_/D vssd1 vssd1 vccd1 vccd1 _18417_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_61_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15629_ _18523_/Q _18487_/Q _15642_/S vssd1 vssd1 vccd1 vccd1 _15629_/X sky130_fd_sc_hd__mux2_1
XFILLER_22_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09150_ _18716_/Q _18715_/Q _18714_/Q vssd1 vssd1 vccd1 vccd1 _09153_/B sky130_fd_sc_hd__or3_4
XFILLER_166_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18348_ _18350_/CLK _18348_/D vssd1 vssd1 vccd1 vccd1 _18348_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_202_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18279_ _18290_/CLK _18279_/D vssd1 vssd1 vccd1 vccd1 _18279_/Q sky130_fd_sc_hd__dfxtp_1
X_09081_ _09083_/A _09081_/B _17833_/Q vssd1 vssd1 vccd1 vccd1 _09082_/A sky130_fd_sc_hd__and3_1
XFILLER_175_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_162_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09983_ _10605_/A _09983_/B _09983_/C vssd1 vssd1 vccd1 vccd1 _13410_/B sky130_fd_sc_hd__and3_1
XFILLER_153_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08934_ _08935_/A vssd1 vssd1 vccd1 vccd1 _08934_/Y sky130_fd_sc_hd__inv_2
XFILLER_229_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_217_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_226_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_213_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_225_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09417_ _18311_/Q _18310_/Q _18309_/Q vssd1 vssd1 vccd1 vccd1 _09418_/D sky130_fd_sc_hd__or3_2
XFILLER_125_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_205_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09348_ _18428_/Q _18427_/Q _18426_/Q vssd1 vssd1 vccd1 vccd1 _09349_/D sky130_fd_sc_hd__or3_4
XFILLER_40_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_200_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_201_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09279_ _18845_/Q _18844_/Q _18843_/Q vssd1 vssd1 vccd1 vccd1 _09282_/B sky130_fd_sc_hd__or3_4
XFILLER_32_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11310_ _11784_/A _11488_/A _11310_/C vssd1 vssd1 vccd1 vccd1 _11491_/A sky130_fd_sc_hd__or3_2
XFILLER_165_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12290_ _12300_/A vssd1 vssd1 vccd1 vccd1 _12327_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_5_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11241_ _11892_/B _11242_/B vssd1 vssd1 vccd1 vccd1 _11243_/B sky130_fd_sc_hd__or2_1
XFILLER_106_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_180_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11172_ _11188_/A vssd1 vssd1 vccd1 vccd1 _11198_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_164_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_212_wb_clk_i clkbuf_5_12_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17793_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_122_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10123_ _10123_/A _10124_/B vssd1 vssd1 vccd1 vccd1 _10129_/B sky130_fd_sc_hd__xnor2_4
X_15980_ _16003_/A _15980_/B vssd1 vssd1 vccd1 vccd1 _15980_/Y sky130_fd_sc_hd__nand2_1
XFILLER_79_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_216_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14931_ _18358_/Q _18322_/Q _14934_/S vssd1 vssd1 vccd1 vccd1 _14931_/X sky130_fd_sc_hd__mux2_1
X_10054_ _09176_/A _09186_/D _10956_/B vssd1 vssd1 vccd1 vccd1 _10054_/X sky130_fd_sc_hd__mux2_1
XFILLER_48_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14862_ _18305_/Q _14861_/B _14861_/Y _14859_/X vssd1 vssd1 vccd1 vccd1 _18305_/D
+ sky130_fd_sc_hd__o211a_1
X_17650_ _17649_/Y _17604_/X _17591_/X vssd1 vssd1 vccd1 vccd1 _17650_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_208_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_217_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16601_ _16599_/B _16598_/X _16599_/Y _16600_/X vssd1 vssd1 vccd1 vccd1 _18719_/D
+ sky130_fd_sc_hd__o211a_1
X_13813_ _18936_/Q _13760_/A _13677_/X _18918_/Q vssd1 vssd1 vccd1 vccd1 _13813_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_4997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17581_ _17581_/A vssd1 vssd1 vccd1 vccd1 _17631_/A sky130_fd_sc_hd__clkbuf_2
X_14793_ _14793_/A _15233_/B _14818_/C vssd1 vssd1 vccd1 vccd1 _14793_/X sky130_fd_sc_hd__or3_1
XFILLER_28_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_217_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16532_ _16555_/A _16678_/B _16568_/C vssd1 vssd1 vccd1 vccd1 _16532_/X sky130_fd_sc_hd__or3_1
XFILLER_216_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13744_ _18321_/Q _13742_/X _13743_/X _18303_/Q vssd1 vssd1 vccd1 vccd1 _13744_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_56_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10956_ _10956_/A _10956_/B vssd1 vssd1 vccd1 vccd1 _10956_/X sky130_fd_sc_hd__or2_1
XFILLER_182_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16463_ _16524_/A vssd1 vssd1 vccd1 vccd1 _16510_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_147_1366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13675_ _18876_/Q _13573_/A _13665_/X _13674_/X vssd1 vssd1 vccd1 vccd1 _13675_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_43_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10887_ _10874_/X _10880_/X _10886_/X _10910_/C vssd1 vssd1 vccd1 vccd1 _10887_/X
+ sky130_fd_sc_hd__o31a_1
XFILLER_32_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15414_ _15417_/B _15412_/X _15413_/Y _15404_/X vssd1 vssd1 vccd1 vccd1 _18436_/D
+ sky130_fd_sc_hd__o211a_1
X_18202_ _18959_/CLK _18202_/D vssd1 vssd1 vccd1 vccd1 _18202_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19182_ _19182_/A _08997_/Y vssd1 vssd1 vccd1 vccd1 io_out[20] sky130_fd_sc_hd__ebufn_8
X_12626_ _12653_/B _12627_/B vssd1 vssd1 vccd1 vccd1 _12628_/A sky130_fd_sc_hd__nand2_1
X_16394_ _16433_/A vssd1 vssd1 vccd1 vccd1 _16452_/B sky130_fd_sc_hd__buf_2
XFILLER_157_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18133_ _18244_/CLK _18133_/D vssd1 vssd1 vccd1 vccd1 _18133_/Q sky130_fd_sc_hd__dfxtp_1
X_15345_ _16853_/A vssd1 vssd1 vccd1 vccd1 _15946_/B sky130_fd_sc_hd__buf_2
XFILLER_8_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_223_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12557_ _12557_/A _12557_/B vssd1 vssd1 vccd1 vccd1 _12557_/Y sky130_fd_sc_hd__nand2_1
XFILLER_184_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18064_ _18072_/CLK _18064_/D vssd1 vssd1 vccd1 vccd1 _18064_/Q sky130_fd_sc_hd__dfxtp_1
X_11508_ _11528_/B _11508_/B _11508_/C vssd1 vssd1 vccd1 vccd1 _11513_/A sky130_fd_sc_hd__and3b_1
X_15276_ _15275_/B _15274_/X _15275_/Y _15264_/X vssd1 vssd1 vccd1 vccd1 _18407_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_129_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_117_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12488_ _12484_/X _12485_/Y _12492_/A _12487_/Y vssd1 vssd1 vccd1 vccd1 _12495_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_156_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17015_ _17015_/A _17449_/B _17028_/C vssd1 vssd1 vccd1 vccd1 _17015_/X sky130_fd_sc_hd__or3_1
X_14227_ _14272_/B vssd1 vssd1 vccd1 vccd1 _14227_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_11439_ _17881_/Q _17880_/Q vssd1 vssd1 vccd1 vccd1 _12323_/B sky130_fd_sc_hd__nand2_1
XFILLER_67_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14158_ _18743_/Q _13546_/X _14154_/X _14157_/X vssd1 vssd1 vccd1 vccd1 _14158_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_4_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13109_ _13142_/A vssd1 vssd1 vccd1 vccd1 _13118_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_140_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14089_ _13434_/C _14073_/X _14080_/X _12027_/B _14088_/X vssd1 vssd1 vccd1 vccd1
+ _14089_/X sky130_fd_sc_hd__a221o_2
X_18966_ _18967_/CLK _18966_/D vssd1 vssd1 vccd1 vccd1 _18966_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_230_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17917_ _18988_/CLK _17917_/D vssd1 vssd1 vccd1 vccd1 _17917_/Q sky130_fd_sc_hd__dfxtp_1
X_18897_ _18899_/CLK _18897_/D vssd1 vssd1 vccd1 vccd1 _18897_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_187_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17848_ _19021_/CLK _17848_/D vssd1 vssd1 vccd1 vccd1 _17848_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_82_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_87_wb_clk_i _18144_/CLK vssd1 vssd1 vccd1 vccd1 _18623_/CLK sky130_fd_sc_hd__clkbuf_16
X_17779_ _18191_/CLK _17779_/D vssd1 vssd1 vccd1 vccd1 _17779_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_19_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_16_wb_clk_i clkbuf_5_5_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18865_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_179_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_228_1176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_1349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_222_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_224_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_223_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09202_ _18587_/Q _18586_/Q _18585_/Q vssd1 vssd1 vccd1 vccd1 _09203_/D sky130_fd_sc_hd__or3_2
XFILLER_22_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09133_ _18824_/Q _18823_/Q _18822_/Q vssd1 vssd1 vccd1 vccd1 _09136_/B sky130_fd_sc_hd__or3_4
XFILLER_163_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09064_ _09064_/A vssd1 vssd1 vccd1 vccd1 _19175_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_120_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_200_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19112__83 vssd1 vssd1 vccd1 vccd1 _19112__83/HI _19220_/A sky130_fd_sc_hd__conb_1
XFILLER_104_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09966_ _12128_/A _09960_/X _09964_/X _10338_/A vssd1 vssd1 vccd1 vccd1 _09966_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_44_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09897_ _09907_/A _09907_/B vssd1 vssd1 vccd1 vccd1 _09924_/A sky130_fd_sc_hd__and2_2
XTAP_4227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_217_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10810_ _09270_/C _09265_/D _10810_/S vssd1 vssd1 vccd1 vccd1 _10811_/B sky130_fd_sc_hd__mux2_1
XFILLER_226_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11790_ _11732_/B _11790_/B vssd1 vssd1 vccd1 vccd1 _11790_/X sky130_fd_sc_hd__and2b_1
XTAP_2869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10741_ _09103_/A _09093_/D _10841_/A vssd1 vssd1 vccd1 vccd1 _10741_/X sky130_fd_sc_hd__mux2_1
XFILLER_25_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_213_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13460_ _17839_/Q _13457_/X _13459_/X vssd1 vssd1 vccd1 vccd1 _13461_/B sky130_fd_sc_hd__a21oi_1
XFILLER_230_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10672_ _10867_/A _10757_/B _10665_/X _10671_/X vssd1 vssd1 vccd1 vccd1 _10672_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_139_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12411_ _17898_/Q _12411_/B vssd1 vssd1 vccd1 vccd1 _12412_/B sky130_fd_sc_hd__and2b_1
X_13391_ _10253_/A _11021_/X _13381_/X _13383_/X vssd1 vssd1 vccd1 vccd1 _18120_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_103_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15130_ _18407_/Q _18371_/Q _15141_/S vssd1 vssd1 vccd1 vccd1 _15130_/X sky130_fd_sc_hd__mux2_1
XFILLER_142_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12342_ _11478_/A _12336_/C _12340_/C _11478_/Y vssd1 vssd1 vccd1 vccd1 _12342_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_126_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15061_ _15061_/A _15061_/B vssd1 vssd1 vccd1 vccd1 _15061_/Y sky130_fd_sc_hd__nand2_1
XFILLER_181_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12273_ _12274_/A _12276_/C _12269_/X _11562_/A _12272_/X vssd1 vssd1 vccd1 vccd1
+ _17867_/D sky130_fd_sc_hd__o221a_1
XFILLER_4_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14012_ _17709_/A _14012_/B vssd1 vssd1 vccd1 vccd1 _14013_/A sky130_fd_sc_hd__or2_1
X_11224_ _11224_/A _17818_/Q _11224_/C vssd1 vssd1 vccd1 vccd1 _11237_/C sky130_fd_sc_hd__and3_1
XFILLER_150_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18820_ _18860_/CLK _18820_/D vssd1 vssd1 vccd1 vccd1 _18820_/Q sky130_fd_sc_hd__dfxtp_4
X_11155_ _11770_/B _17813_/Q _12285_/A vssd1 vssd1 vccd1 vccd1 _11156_/A sky130_fd_sc_hd__mux2_1
XFILLER_96_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10106_ _09694_/A _10101_/X _10105_/X _10044_/A vssd1 vssd1 vccd1 vccd1 _10106_/X
+ sky130_fd_sc_hd__o211a_1
X_18751_ _18752_/CLK _18751_/D vssd1 vssd1 vccd1 vccd1 _18751_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_62_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15963_ _18603_/Q _18567_/Q _15963_/S vssd1 vssd1 vccd1 vccd1 _15963_/X sky130_fd_sc_hd__mux2_1
XTAP_5440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11086_ _12023_/A vssd1 vssd1 vccd1 vccd1 _11313_/B sky130_fd_sc_hd__clkbuf_2
XTAP_5451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17702_ _18988_/Q _17701_/Y _17705_/S vssd1 vssd1 vccd1 vccd1 _17703_/A sky130_fd_sc_hd__mux2_1
X_14914_ _14913_/B _14912_/X _14913_/Y _14902_/X vssd1 vssd1 vccd1 vccd1 _18317_/D
+ sky130_fd_sc_hd__o211a_1
X_10037_ _09165_/A _09160_/C _09170_/D _10308_/A _10036_/X _09986_/A vssd1 vssd1 vccd1
+ vccd1 _10037_/X sky130_fd_sc_hd__mux4_1
XFILLER_114_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18682_ _18682_/CLK _18682_/D vssd1 vssd1 vccd1 vccd1 _18682_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_5484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15894_ _15921_/A _16043_/B _15894_/C vssd1 vssd1 vccd1 vccd1 _15894_/X sky130_fd_sc_hd__or3_1
XTAP_5495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_224_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17633_ _17638_/A _17633_/B vssd1 vssd1 vccd1 vccd1 _17634_/A sky130_fd_sc_hd__and2_1
X_14845_ _18337_/Q _18301_/Q _14848_/S vssd1 vssd1 vccd1 vccd1 _14845_/X sky130_fd_sc_hd__mux2_1
XFILLER_36_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_217_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14776_ _18283_/Q _14777_/B _14775_/Y _14758_/X vssd1 vssd1 vccd1 vccd1 _18283_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_16_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17564_ _17564_/A _17564_/B vssd1 vssd1 vccd1 vccd1 _17565_/A sky130_fd_sc_hd__and2_1
XFILLER_223_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11988_ _11988_/A _12007_/B _11988_/C vssd1 vssd1 vccd1 vccd1 _13434_/C sky130_fd_sc_hd__nor3_4
XFILLER_90_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16515_ _16807_/A _16652_/C vssd1 vssd1 vccd1 vccd1 _16525_/B sky130_fd_sc_hd__nor2_1
X_13727_ _18261_/Q _13615_/A _13722_/X _13726_/X vssd1 vssd1 vccd1 vccd1 _13727_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_108_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10939_ _10939_/A _10939_/B _10939_/C vssd1 vssd1 vccd1 vccd1 _10939_/X sky130_fd_sc_hd__or3_1
XFILLER_205_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17495_ _18973_/Q _18937_/Q _17495_/S vssd1 vssd1 vccd1 vccd1 _17495_/X sky130_fd_sc_hd__mux2_1
XFILLER_189_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19234_ _19234_/A _08938_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[34] sky130_fd_sc_hd__ebufn_8
XFILLER_220_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16446_ _18718_/Q _18682_/Q _16449_/S vssd1 vssd1 vccd1 vccd1 _16446_/X sky130_fd_sc_hd__mux2_1
X_13658_ _18954_/Q _13642_/A _13513_/A _18960_/Q vssd1 vssd1 vccd1 vccd1 _13658_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_231_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_220_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12609_ _12637_/B _12609_/B vssd1 vssd1 vccd1 vccd1 _12610_/B sky130_fd_sc_hd__and2_1
X_19165_ _19165_/A _09028_/Y vssd1 vssd1 vccd1 vccd1 io_out[3] sky130_fd_sc_hd__ebufn_8
X_16377_ _18664_/Q _16378_/B _16373_/Y _16376_/X vssd1 vssd1 vccd1 vccd1 _18664_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_185_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13589_ _18720_/Q _13856_/A _13588_/X _18711_/Q vssd1 vssd1 vccd1 vccd1 _13589_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_34_1366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15328_ _15370_/A vssd1 vssd1 vccd1 vccd1 _15393_/B sky130_fd_sc_hd__buf_2
XFILLER_173_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18116_ _18125_/CLK _18116_/D vssd1 vssd1 vccd1 vccd1 _18116_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_219_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_134_wb_clk_i clkbuf_5_27_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18374_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_117_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15259_ _18439_/Q _18403_/Q _15267_/S vssd1 vssd1 vccd1 vccd1 _15259_/X sky130_fd_sc_hd__mux2_1
XFILLER_144_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18047_ _18052_/CLK _18047_/D vssd1 vssd1 vccd1 vccd1 _18047_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_160_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_125_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09820_ _12131_/A _12133_/A vssd1 vssd1 vccd1 vccd1 _09983_/B sky130_fd_sc_hd__and2b_1
XFILLER_99_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_193_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09751_ _09751_/A _09751_/B vssd1 vssd1 vccd1 vccd1 _09816_/A sky130_fd_sc_hd__or2_1
XFILLER_98_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18949_ _18950_/CLK _18949_/D vssd1 vssd1 vccd1 vccd1 _18949_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_228_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09682_ _09682_/A vssd1 vssd1 vccd1 vccd1 _10085_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_55_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_228_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_215_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09116_ _18743_/Q _18742_/Q _18741_/Q vssd1 vssd1 vccd1 vccd1 _09119_/B sky130_fd_sc_hd__or3_4
XFILLER_136_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09047_ _09053_/A vssd1 vssd1 vccd1 vccd1 _09052_/A sky130_fd_sc_hd__buf_12
XFILLER_89_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09949_ _09397_/A _09392_/D _12124_/A vssd1 vssd1 vccd1 vccd1 _09949_/X sky130_fd_sc_hd__mux2_1
XFILLER_213_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12960_ _12961_/A _12961_/B vssd1 vssd1 vccd1 vccd1 _12960_/X sky130_fd_sc_hd__or2_1
XFILLER_58_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XINSDIODE2_30 _10990_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_180_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_41 _10940_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_52 _10772_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_63 _12318_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11911_ _10264_/A _10264_/B _11910_/Y vssd1 vssd1 vccd1 vccd1 _11919_/A sky130_fd_sc_hd__a21o_1
XINSDIODE2_74 _13576_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12891_ _17960_/Q _12890_/B _12854_/X vssd1 vssd1 vccd1 vccd1 _12892_/B sky130_fd_sc_hd__o21ai_1
XFILLER_79_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XINSDIODE2_85 _13621_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_96 _13739_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14630_ _18249_/Q _14635_/B _14628_/X _14629_/X vssd1 vssd1 vccd1 vccd1 _18249_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_3378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11842_ _11842_/A _11842_/B _11842_/C vssd1 vssd1 vccd1 vccd1 _11845_/B sky130_fd_sc_hd__or3_1
XFILLER_57_1300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14561_ _14668_/A vssd1 vssd1 vccd1 vccd1 _14561_/X sky130_fd_sc_hd__clkbuf_2
XTAP_1943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11773_ _11769_/X _11772_/X _11763_/X _11765_/X vssd1 vssd1 vccd1 vccd1 _11773_/X
+ sky130_fd_sc_hd__o2bb2a_1
XTAP_1954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16300_ _16305_/B _16298_/X _16299_/X _16295_/X vssd1 vssd1 vccd1 vccd1 _18645_/D
+ sky130_fd_sc_hd__o211a_1
X_13512_ _13734_/A vssd1 vssd1 vccd1 vccd1 _13513_/A sky130_fd_sc_hd__clkbuf_4
XTAP_1976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10724_ _10664_/A _10720_/X _10723_/X _10818_/A vssd1 vssd1 vccd1 vccd1 _10724_/X
+ sky130_fd_sc_hd__a211o_1
XTAP_1987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17280_ _17370_/A vssd1 vssd1 vccd1 vccd1 _17298_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_213_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14492_ _14492_/A vssd1 vssd1 vccd1 vccd1 _18220_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16231_ _18629_/Q _16229_/B _16229_/Y _16230_/X vssd1 vssd1 vccd1 vccd1 _18629_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_13_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13443_ _13443_/A _13452_/B vssd1 vssd1 vccd1 vccd1 _13443_/Y sky130_fd_sc_hd__nor2_1
XFILLER_13_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10655_ _10818_/B vssd1 vssd1 vccd1 vccd1 _10757_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_186_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16162_ _16252_/A vssd1 vssd1 vccd1 vccd1 _16162_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_155_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13374_ _18110_/Q _13389_/B vssd1 vssd1 vccd1 vccd1 _13374_/Y sky130_fd_sc_hd__nand2_1
XFILLER_154_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10586_ _09314_/A _09319_/B _09314_/D _09314_/C _09688_/A _09682_/A vssd1 vssd1 vccd1
+ vccd1 _10586_/X sky130_fd_sc_hd__mux4_1
XFILLER_186_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15113_ _15118_/B _15110_/X _15112_/X _15103_/X vssd1 vssd1 vccd1 vccd1 _18366_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_127_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12325_ _13153_/A _12325_/B vssd1 vssd1 vccd1 vccd1 _17881_/D sky130_fd_sc_hd__nor2_1
X_16093_ _16096_/B _16091_/X _16092_/Y _16074_/X vssd1 vssd1 vccd1 vccd1 _18598_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_114_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15044_ _18385_/Q _18349_/Q _15052_/S vssd1 vssd1 vccd1 vccd1 _15044_/X sky130_fd_sc_hd__mux2_1
XFILLER_138_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12256_ _17863_/Q _12253_/Y _12276_/C _12219_/X vssd1 vssd1 vccd1 vccd1 _17863_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_170_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_2_1_0_wb_clk_i clkbuf_2_1_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_2_1_1_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_2
X_11207_ _11207_/A vssd1 vssd1 vccd1 vccd1 _17813_/D sky130_fd_sc_hd__clkbuf_1
X_12187_ _18106_/Q _18990_/Q _18991_/Q _12401_/B vssd1 vssd1 vccd1 vccd1 _12444_/B
+ sky130_fd_sc_hd__or4_4
XFILLER_123_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_218_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18803_ _18806_/CLK _18803_/D vssd1 vssd1 vccd1 vccd1 _18803_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_150_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11138_ _11138_/A vssd1 vssd1 vccd1 vccd1 _17800_/D sky130_fd_sc_hd__clkbuf_1
X_16995_ _17032_/A _16998_/B vssd1 vssd1 vccd1 vccd1 _16995_/Y sky130_fd_sc_hd__nand2_1
XFILLER_23_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18734_ _18765_/CLK _18734_/D vssd1 vssd1 vccd1 vccd1 _18734_/Q sky130_fd_sc_hd__dfxtp_1
X_15946_ _15984_/A _15946_/B _15964_/C vssd1 vssd1 vccd1 vccd1 _15946_/X sky130_fd_sc_hd__or3_1
XTAP_5270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11069_ _11368_/B vssd1 vssd1 vccd1 vccd1 _13442_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_110_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_209_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18665_ _18696_/CLK _18665_/D vssd1 vssd1 vccd1 vccd1 _18665_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_48_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15877_ _15876_/B _15875_/X _15876_/Y _15861_/X vssd1 vssd1 vccd1 vccd1 _18548_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_4580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_225_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17616_ _17687_/B _17663_/A vssd1 vssd1 vccd1 vccd1 _17616_/Y sky130_fd_sc_hd__nor2_1
XFILLER_92_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14828_ _14827_/B _14825_/X _14827_/Y _14819_/X vssd1 vssd1 vccd1 vccd1 _18296_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_52_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18596_ _18608_/CLK _18596_/D vssd1 vssd1 vccd1 vccd1 _18596_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_92_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_225_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17547_ _17547_/A vssd1 vssd1 vccd1 vccd1 _17547_/X sky130_fd_sc_hd__clkbuf_2
X_14759_ _14767_/B _14756_/X _14757_/X _14758_/X vssd1 vssd1 vccd1 vccd1 _18279_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_44_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_225_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_220_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17478_ _17497_/A vssd1 vssd1 vccd1 vccd1 _17478_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_149_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19217_ _19217_/A _08970_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[17] sky130_fd_sc_hd__ebufn_8
X_16429_ _16450_/A _16429_/B vssd1 vssd1 vccd1 vccd1 _16429_/Y sky130_fd_sc_hd__nand2_1
XFILLER_34_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19148_ _19148_/A _09040_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[18] sky130_fd_sc_hd__ebufn_8
XFILLER_34_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_191_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_195_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09803_ _09743_/A _10675_/A _09742_/A vssd1 vssd1 vccd1 vccd1 _09803_/X sky130_fd_sc_hd__a21o_1
XFILLER_101_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_1240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09734_ _19027_/Q _17979_/Q vssd1 vssd1 vccd1 vccd1 _10116_/B sky130_fd_sc_hd__xor2_4
XFILLER_28_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_31_wb_clk_i clkbuf_5_7_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18950_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_80_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09665_ _09665_/A _09665_/B vssd1 vssd1 vccd1 vccd1 _09665_/X sky130_fd_sc_hd__or2_1
XFILLER_216_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09596_ _09725_/B _09725_/A vssd1 vssd1 vccd1 vccd1 _09596_/X sky130_fd_sc_hd__and2b_1
XFILLER_199_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_211_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_210_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10440_ _10440_/A _10440_/B vssd1 vssd1 vccd1 vccd1 _10441_/B sky130_fd_sc_hd__and2_1
XFILLER_52_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10371_ _09889_/A _10367_/X _10370_/X _09981_/A vssd1 vssd1 vccd1 vccd1 _10371_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_164_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12110_ _09822_/A _09844_/A _09843_/B _12109_/X vssd1 vssd1 vccd1 vccd1 _12118_/A
+ sky130_fd_sc_hd__a31o_1
XFILLER_108_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13090_ _18006_/Q _14377_/A vssd1 vssd1 vccd1 vccd1 _13091_/A sky130_fd_sc_hd__or2_1
XFILLER_123_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12041_ _12041_/A _12041_/B _12041_/C vssd1 vssd1 vccd1 vccd1 _12042_/B sky130_fd_sc_hd__nor3_4
XFILLER_104_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_215_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15800_ _15806_/B _15798_/X _15799_/X _15783_/X vssd1 vssd1 vccd1 vccd1 _18528_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_213_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13992_ _12019_/B _13984_/X _13991_/X _12055_/B vssd1 vssd1 vccd1 vccd1 _13992_/X
+ sky130_fd_sc_hd__a22o_2
X_16780_ _16780_/A vssd1 vssd1 vccd1 vccd1 _16871_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_19_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_219_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15731_ _15730_/B _15729_/X _15730_/Y _15720_/X vssd1 vssd1 vccd1 vccd1 _18512_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_20_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12943_ _17995_/Q _12955_/A _12933_/A _12941_/Y _13368_/A vssd1 vssd1 vccd1 vccd1
+ _12944_/B sky130_fd_sc_hd__a32o_1
XTAP_3120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_219_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18450_ _18467_/CLK _18450_/D vssd1 vssd1 vccd1 vccd1 _18450_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_34_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15662_ _15720_/A vssd1 vssd1 vccd1 vccd1 _15662_/X sky130_fd_sc_hd__clkbuf_2
X_12874_ _12874_/A vssd1 vssd1 vccd1 vccd1 _12874_/X sky130_fd_sc_hd__clkbuf_2
XTAP_2430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17401_ _17408_/B _17398_/X _17399_/X _17400_/X vssd1 vssd1 vccd1 vccd1 _18912_/D
+ sky130_fd_sc_hd__o211a_1
X_14613_ _14608_/X _14612_/A _18246_/Q vssd1 vssd1 vccd1 vccd1 _14613_/Y sky130_fd_sc_hd__o21bai_1
X_11825_ _11826_/A _11826_/B _11826_/C vssd1 vssd1 vccd1 vccd1 _11825_/Y sky130_fd_sc_hd__o21ai_1
X_18381_ _18392_/CLK _18381_/D vssd1 vssd1 vccd1 vccd1 _18381_/Q sky130_fd_sc_hd__dfxtp_2
X_15593_ _18515_/Q _18479_/Q _15604_/S vssd1 vssd1 vccd1 vccd1 _15593_/X sky130_fd_sc_hd__mux2_1
XFILLER_33_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14544_ _17544_/A vssd1 vssd1 vccd1 vccd1 _14606_/A sky130_fd_sc_hd__clkbuf_2
XTAP_1773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17332_ _17376_/A _17473_/B _17376_/C vssd1 vssd1 vccd1 vccd1 _17332_/X sky130_fd_sc_hd__or3_1
XFILLER_14_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11756_ _11767_/C _11753_/X _11756_/S vssd1 vssd1 vccd1 vccd1 _11797_/A sky130_fd_sc_hd__mux2_1
XTAP_1784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_186_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_197_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10707_ _10843_/B _12101_/A vssd1 vssd1 vccd1 vccd1 _10707_/Y sky130_fd_sc_hd__nor2_1
XFILLER_41_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14475_ _14475_/A vssd1 vssd1 vccd1 vccd1 _18212_/D sky130_fd_sc_hd__clkbuf_1
X_17263_ _17275_/A _17263_/B vssd1 vssd1 vccd1 vccd1 _17263_/Y sky130_fd_sc_hd__nand2_1
X_11687_ _17852_/Q _11703_/A vssd1 vssd1 vccd1 vccd1 _11687_/Y sky130_fd_sc_hd__nor2_1
XFILLER_70_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19002_ _19004_/CLK _19002_/D vssd1 vssd1 vccd1 vccd1 _19002_/Q sky130_fd_sc_hd__dfxtp_1
X_16214_ _16217_/B _16211_/X _16213_/Y _16209_/X vssd1 vssd1 vccd1 vccd1 _18625_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_174_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13426_ _13426_/A _13426_/B vssd1 vssd1 vccd1 vccd1 _13426_/Y sky130_fd_sc_hd__xnor2_4
X_10638_ _10667_/A vssd1 vssd1 vccd1 vccd1 _10766_/A sky130_fd_sc_hd__clkbuf_2
X_17194_ _17200_/B _17192_/X _17193_/X _17181_/X vssd1 vssd1 vccd1 vccd1 _18861_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_155_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16145_ _18647_/Q _18611_/Q _16145_/S vssd1 vssd1 vccd1 vccd1 _16145_/X sky130_fd_sc_hd__mux2_1
XFILLER_10_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13357_ _18131_/Q _13357_/B vssd1 vssd1 vccd1 vccd1 _14422_/A sky130_fd_sc_hd__nand2_4
X_10569_ _10569_/A _10575_/B vssd1 vssd1 vccd1 vccd1 _10569_/X sky130_fd_sc_hd__or2_1
XFILLER_155_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12308_ _11323_/X _12292_/B _12329_/C _12307_/Y _11891_/X vssd1 vssd1 vccd1 vccd1
+ _17877_/D sky130_fd_sc_hd__a2111oi_1
XFILLER_5_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16076_ _18631_/Q _18595_/Q _16091_/S vssd1 vssd1 vccd1 vccd1 _16076_/X sky130_fd_sc_hd__mux2_1
X_13288_ _18021_/Q _18020_/Q _18023_/Q _18022_/Q vssd1 vssd1 vccd1 vccd1 _13291_/B
+ sky130_fd_sc_hd__or4_1
XFILLER_170_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15027_ _15025_/B _15024_/X _15025_/Y _15026_/X vssd1 vssd1 vccd1 vccd1 _18344_/D
+ sky130_fd_sc_hd__o211a_1
X_12239_ _17859_/Q _17556_/A _12239_/C vssd1 vssd1 vccd1 vccd1 _12240_/A sky130_fd_sc_hd__and3_1
XFILLER_155_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_1268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_231_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16978_ _17107_/B vssd1 vssd1 vccd1 vccd1 _16978_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_83_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput4 io_in[26] vssd1 vssd1 vccd1 vccd1 input4/X sky130_fd_sc_hd__clkbuf_1
XFILLER_49_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18717_ _18722_/CLK _18717_/D vssd1 vssd1 vccd1 vccd1 _18717_/Q sky130_fd_sc_hd__dfxtp_4
X_15929_ _15928_/B _15927_/X _15928_/Y _15925_/X vssd1 vssd1 vccd1 vccd1 _18560_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_209_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09450_ _09450_/A _09450_/B vssd1 vssd1 vccd1 vccd1 _09450_/Y sky130_fd_sc_hd__nor2_1
XFILLER_224_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18648_ _18668_/CLK _18648_/D vssd1 vssd1 vccd1 vccd1 _18648_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_225_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_224_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09381_ _09381_/A _09381_/B _09381_/C _09381_/D vssd1 vssd1 vccd1 vccd1 _09387_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_149_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18579_ _18582_/CLK _18579_/D vssd1 vssd1 vccd1 vccd1 _18579_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_75_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_221_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_220_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_220_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_220_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_105_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_1335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_216_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09717_ _10065_/A vssd1 vssd1 vccd1 vccd1 _10944_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_56_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09648_ _09664_/A _09684_/B vssd1 vssd1 vccd1 vccd1 _09704_/A sky130_fd_sc_hd__nor2_1
XTAP_1003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_216_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09579_ _17980_/Q vssd1 vssd1 vccd1 vccd1 _10705_/A sky130_fd_sc_hd__buf_4
XTAP_1047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11610_ _11603_/Y _11608_/X _11609_/X vssd1 vssd1 vccd1 vccd1 _11610_/Y sky130_fd_sc_hd__a21oi_1
XTAP_1069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12590_ _12590_/A _12590_/B vssd1 vssd1 vccd1 vccd1 _12590_/Y sky130_fd_sc_hd__nand2_1
XFILLER_143_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_1366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11541_ _11541_/A _11541_/B vssd1 vssd1 vccd1 vccd1 _11921_/B sky130_fd_sc_hd__nand2_1
XFILLER_54_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_184_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_168_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14260_ _14260_/A _14260_/B vssd1 vssd1 vccd1 vccd1 _14260_/Y sky130_fd_sc_hd__nand2_1
XFILLER_156_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11472_ _11472_/A _12337_/S vssd1 vssd1 vccd1 vccd1 _11478_/B sky130_fd_sc_hd__nor2_1
XFILLER_184_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13211_ _13467_/A input5/X vssd1 vssd1 vccd1 vccd1 _18061_/D sky130_fd_sc_hd__nor2_1
XFILLER_52_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10423_ _14307_/A _12047_/A vssd1 vssd1 vccd1 vccd1 _10533_/B sky130_fd_sc_hd__or2_2
X_14191_ _18207_/Q vssd1 vssd1 vccd1 vccd1 _14233_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_136_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13142_ _13142_/A vssd1 vssd1 vccd1 vccd1 _13151_/A sky130_fd_sc_hd__clkbuf_1
X_10354_ _09993_/A _09153_/B _09148_/A _09143_/D _10274_/S _09905_/X vssd1 vssd1 vccd1
+ vccd1 _10354_/X sky130_fd_sc_hd__mux4_2
XFILLER_191_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17950_ _17954_/CLK _17950_/D vssd1 vssd1 vccd1 vccd1 _17950_/Q sky130_fd_sc_hd__dfxtp_1
X_13073_ _17747_/A vssd1 vssd1 vccd1 vccd1 _14533_/A sky130_fd_sc_hd__clkbuf_4
X_10285_ _09219_/B _09214_/B _10285_/S vssd1 vssd1 vccd1 vccd1 _10285_/X sky130_fd_sc_hd__mux2_1
XFILLER_2_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_219_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16901_ _17228_/A vssd1 vssd1 vccd1 vccd1 _17168_/A sky130_fd_sc_hd__clkbuf_2
X_12024_ _11974_/B _11591_/B _12023_/Y _12026_/B _12007_/B vssd1 vssd1 vccd1 vccd1
+ _12027_/A sky130_fd_sc_hd__o311a_4
XFILLER_78_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_215_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17881_ _17883_/CLK _17881_/D vssd1 vssd1 vccd1 vccd1 _17881_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_215_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16832_ _16832_/A vssd1 vssd1 vccd1 vccd1 _16884_/A sky130_fd_sc_hd__buf_2
XFILLER_93_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19073__44 vssd1 vssd1 vccd1 vccd1 _19073__44/HI _19167_/A sky130_fd_sc_hd__conb_1
XFILLER_76_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_219_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16763_ _16828_/A vssd1 vssd1 vccd1 vccd1 _16813_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_20_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13975_ _18298_/Q _13738_/X _13973_/X _13974_/X vssd1 vssd1 vccd1 vccd1 _13975_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_24_1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18502_ _18532_/CLK _18502_/D vssd1 vssd1 vccd1 vccd1 _18502_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_47_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15714_ _18544_/Q _18508_/Q _15714_/S vssd1 vssd1 vccd1 vccd1 _15714_/X sky130_fd_sc_hd__mux2_1
XFILLER_94_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_206_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12926_ _12926_/A _13041_/A vssd1 vssd1 vccd1 vccd1 _12931_/A sky130_fd_sc_hd__nor2_1
XFILLER_185_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16694_ _18778_/Q _18742_/Q _16694_/S vssd1 vssd1 vccd1 vccd1 _16694_/X sky130_fd_sc_hd__mux2_1
XFILLER_18_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18433_ _18434_/CLK _18433_/D vssd1 vssd1 vccd1 vccd1 _18433_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_146_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15645_ _15691_/A _15651_/B vssd1 vssd1 vccd1 vccd1 _15645_/Y sky130_fd_sc_hd__nand2_1
XTAP_2260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12857_ _17949_/Q _17950_/Q _12857_/C vssd1 vssd1 vccd1 vccd1 _12865_/C sky130_fd_sc_hd__and3_1
XTAP_2271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_226_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18364_ _18392_/CLK _18364_/D vssd1 vssd1 vccd1 vccd1 _18364_/Q sky130_fd_sc_hd__dfxtp_2
X_11808_ _11812_/B _11808_/B _11808_/C _11807_/X vssd1 vssd1 vccd1 vccd1 _11869_/B
+ sky130_fd_sc_hd__or4b_4
XFILLER_199_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15576_ _15583_/B _15573_/X _15574_/X _15575_/X vssd1 vssd1 vccd1 vccd1 _18474_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_1570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12788_ _13080_/A _13082_/A vssd1 vssd1 vccd1 vccd1 _12788_/Y sky130_fd_sc_hd__nor2_1
XFILLER_187_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17315_ _17314_/B _17313_/X _17314_/Y _17304_/X vssd1 vssd1 vccd1 vccd1 _18890_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_230_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14527_ _14598_/A vssd1 vssd1 vccd1 vccd1 _14690_/B sky130_fd_sc_hd__buf_2
XFILLER_14_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11739_ _11727_/A _11767_/C _11760_/B _11747_/A vssd1 vssd1 vccd1 vccd1 _11740_/C
+ sky130_fd_sc_hd__o22a_1
XFILLER_159_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18295_ _18308_/CLK _18295_/D vssd1 vssd1 vccd1 vccd1 _18295_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_222_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17246_ _17252_/B _17244_/X _17245_/X _17241_/X vssd1 vssd1 vccd1 vccd1 _18873_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_186_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14458_ _14458_/A vssd1 vssd1 vccd1 vccd1 _18205_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_190_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_179_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_122_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13409_ _14299_/A vssd1 vssd1 vccd1 vccd1 _13409_/X sky130_fd_sc_hd__clkbuf_4
X_14389_ _17661_/A vssd1 vssd1 vccd1 vccd1 _17640_/A sky130_fd_sc_hd__clkbuf_2
X_17177_ _17210_/A _17180_/B vssd1 vssd1 vccd1 vccd1 _17177_/Y sky130_fd_sc_hd__nand2_1
XFILLER_31_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16128_ _16181_/A _16128_/B _16181_/C vssd1 vssd1 vccd1 vccd1 _16128_/X sky130_fd_sc_hd__or3_1
XFILLER_155_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08950_ _08954_/A vssd1 vssd1 vccd1 vccd1 _08950_/Y sky130_fd_sc_hd__inv_2
X_16059_ _16205_/B vssd1 vssd1 vccd1 vccd1 _16115_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_115_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_217_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_1240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09502_ _18200_/Q _09502_/B vssd1 vssd1 vccd1 vccd1 _09503_/B sky130_fd_sc_hd__or2_1
XFILLER_112_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09433_ _09435_/B _09482_/A vssd1 vssd1 vccd1 vccd1 _09434_/A sky130_fd_sc_hd__and2b_1
XFILLER_164_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09364_ _18287_/Q _18286_/Q _18285_/Q vssd1 vssd1 vccd1 vccd1 _09365_/D sky130_fd_sc_hd__or3_4
XFILLER_24_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_197_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_205_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09295_ _18518_/Q _18517_/Q _18516_/Q vssd1 vssd1 vccd1 vccd1 _10569_/A sky130_fd_sc_hd__or3_4
XFILLER_21_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_192_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10070_ _10033_/A _10070_/B vssd1 vssd1 vccd1 vccd1 _10966_/B sky130_fd_sc_hd__and2b_4
XTAP_5814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_1176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13760_ _13760_/A vssd1 vssd1 vccd1 vccd1 _13847_/A sky130_fd_sc_hd__buf_6
XFILLER_21_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10972_ _14507_/A _13417_/B vssd1 vssd1 vccd1 vccd1 _13412_/C sky130_fd_sc_hd__and2_1
XFILLER_216_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_231_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_204_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12711_ _17938_/Q _12707_/X _12710_/Y vssd1 vssd1 vccd1 vccd1 _17938_/D sky130_fd_sc_hd__a21o_1
X_13691_ _18621_/Q _13657_/A _13689_/X _13690_/X vssd1 vssd1 vccd1 vccd1 _13691_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_188_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_203_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_231_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15430_ _18476_/Q _18440_/Q _15435_/S vssd1 vssd1 vccd1 vccd1 _15430_/X sky130_fd_sc_hd__mux2_1
X_12642_ _17928_/Q _12635_/X _12640_/Y _12641_/X _12621_/X vssd1 vssd1 vccd1 vccd1
+ _17928_/D sky130_fd_sc_hd__a221o_1
XFILLER_93_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_93_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_231_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15361_ _18460_/Q _18424_/Q _15388_/S vssd1 vssd1 vccd1 vccd1 _15361_/X sky130_fd_sc_hd__mux2_1
X_12573_ _12573_/A vssd1 vssd1 vccd1 vccd1 _12575_/A sky130_fd_sc_hd__inv_2
XFILLER_178_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_197_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17100_ _17164_/A vssd1 vssd1 vccd1 vccd1 _17152_/A sky130_fd_sc_hd__buf_2
XFILLER_12_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11524_ _11513_/A _11520_/X _11523_/X _11526_/B vssd1 vssd1 vccd1 vccd1 _11524_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_11_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14312_ _14355_/B _14321_/A vssd1 vssd1 vccd1 vccd1 _14312_/X sky130_fd_sc_hd__or2_1
X_15292_ _15292_/A _15451_/C vssd1 vssd1 vccd1 vccd1 _15303_/B sky130_fd_sc_hd__nor2_2
X_18080_ _18087_/CLK _18080_/D vssd1 vssd1 vccd1 vccd1 _18080_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_178_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17031_ _18856_/Q _18820_/Q _17055_/S vssd1 vssd1 vccd1 vccd1 _17031_/X sky130_fd_sc_hd__mux2_1
X_14243_ _14299_/A vssd1 vssd1 vccd1 vccd1 _14243_/X sky130_fd_sc_hd__clkbuf_2
X_11455_ _11374_/B _13429_/A _11455_/C _11455_/D vssd1 vssd1 vccd1 vccd1 _11455_/X
+ sky130_fd_sc_hd__and4b_1
XFILLER_194_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10406_ _10605_/A vssd1 vssd1 vccd1 vccd1 _10406_/Y sky130_fd_sc_hd__inv_2
X_14174_ _18626_/Q _13612_/X _14027_/X _18617_/Q _14173_/X vssd1 vssd1 vccd1 vccd1
+ _14174_/X sky130_fd_sc_hd__a221o_1
X_11386_ _11331_/X _11385_/X _11346_/Y vssd1 vssd1 vccd1 vccd1 _11386_/X sky130_fd_sc_hd__o21a_1
XFILLER_124_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13125_ _13129_/A _18023_/Q vssd1 vssd1 vccd1 vccd1 _13126_/A sky130_fd_sc_hd__and2_1
XFILLER_113_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10337_ _09143_/C _09148_/B _09153_/D _09148_/D _09909_/X _12121_/A vssd1 vssd1 vccd1
+ vccd1 _10338_/B sky130_fd_sc_hd__mux4_2
X_18982_ _18986_/CLK _18982_/D vssd1 vssd1 vccd1 vccd1 _18982_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_97_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13056_ _13054_/Y _13055_/X _13066_/C vssd1 vssd1 vccd1 vccd1 _13056_/X sky130_fd_sc_hd__a21o_1
X_17933_ _17933_/CLK _17933_/D vssd1 vssd1 vccd1 vccd1 _17933_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_26_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10268_ _10513_/A vssd1 vssd1 vccd1 vccd1 _10918_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_191_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12007_ _12007_/A _12007_/B vssd1 vssd1 vccd1 vccd1 _12007_/Y sky130_fd_sc_hd__nand2_1
XFILLER_6_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17864_ _17864_/CLK _17864_/D vssd1 vssd1 vccd1 vccd1 _17864_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_113_1216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10199_ _10197_/A _10197_/B _10202_/A vssd1 vssd1 vccd1 vccd1 _10246_/B sky130_fd_sc_hd__o21ba_1
Xclkbuf_leaf_159_wb_clk_i _18114_/CLK vssd1 vssd1 vccd1 vccd1 _19027_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_93_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16815_ _16815_/A _16815_/B vssd1 vssd1 vccd1 vccd1 _16815_/Y sky130_fd_sc_hd__nand2_1
X_17795_ _17806_/CLK _17795_/D vssd1 vssd1 vccd1 vccd1 _17795_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_94_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_219_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16746_ _16766_/A vssd1 vssd1 vccd1 vccd1 _16762_/S sky130_fd_sc_hd__clkbuf_2
X_13958_ _18631_/Q _13719_/X _13721_/X _18655_/Q vssd1 vssd1 vccd1 vccd1 _13958_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_4_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_228_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12909_ _17966_/Q _12908_/B _12854_/X vssd1 vssd1 vccd1 vccd1 _12910_/B sky130_fd_sc_hd__o21ai_1
XFILLER_185_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16677_ _18774_/Q _18738_/Q _16694_/S vssd1 vssd1 vccd1 vccd1 _16677_/X sky130_fd_sc_hd__mux2_1
X_13889_ _18958_/Q _13651_/X _13885_/X _13888_/X vssd1 vssd1 vccd1 vccd1 _13889_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_228_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18416_ _18416_/CLK _18416_/D vssd1 vssd1 vccd1 vccd1 _18416_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_34_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15628_ _15633_/B _15624_/X _15627_/X _15616_/X vssd1 vssd1 vccd1 vccd1 _18486_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_179_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_222_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_222_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18347_ _18367_/CLK _18347_/D vssd1 vssd1 vccd1 vccd1 _18347_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_21_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_226_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15559_ _15558_/B _15557_/X _15558_/Y _15555_/X vssd1 vssd1 vccd1 vccd1 _18470_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_187_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09080_ _09080_/A vssd1 vssd1 vccd1 vccd1 _19186_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_174_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18278_ _18278_/CLK _18278_/D vssd1 vssd1 vccd1 vccd1 _18278_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_200_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17229_ _17468_/A vssd1 vssd1 vccd1 vccd1 _17275_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_174_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_128_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09982_ _09889_/X _09932_/X _09978_/X _09981_/X vssd1 vssd1 vccd1 vccd1 _09983_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_116_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08933_ _08935_/A vssd1 vssd1 vccd1 vccd1 _08933_/Y sky130_fd_sc_hd__inv_2
XFILLER_103_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_226_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_225_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09416_ _18335_/Q _18334_/Q _18333_/Q vssd1 vssd1 vccd1 vccd1 _09418_/C sky130_fd_sc_hd__or3_1
XFILLER_13_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_179_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09347_ _18419_/Q _18418_/Q _18417_/Q vssd1 vssd1 vccd1 vccd1 _10391_/A sky130_fd_sc_hd__or3_4
XFILLER_205_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09278_ _18866_/Q _18865_/Q _18864_/Q vssd1 vssd1 vccd1 vccd1 _09282_/A sky130_fd_sc_hd__or3_4
XFILLER_138_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11240_ _11240_/A vssd1 vssd1 vccd1 vccd1 _17822_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_153_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11171_ _11209_/A _17813_/Q _11169_/X _17661_/A vssd1 vssd1 vccd1 vccd1 _11188_/A
+ sky130_fd_sc_hd__o31a_1
XFILLER_122_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10122_ _10122_/A _10122_/B vssd1 vssd1 vccd1 vccd1 _10124_/B sky130_fd_sc_hd__xnor2_4
XFILLER_164_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_216_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14930_ _14935_/B _14927_/X _14929_/X _14922_/X vssd1 vssd1 vccd1 vccd1 _18321_/D
+ sky130_fd_sc_hd__o211a_1
X_10053_ _10053_/A _10053_/B vssd1 vssd1 vccd1 vccd1 _10053_/X sky130_fd_sc_hd__or2_1
XTAP_5644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14861_ _14875_/A _14861_/B vssd1 vssd1 vccd1 vccd1 _14861_/Y sky130_fd_sc_hd__nand2_1
XTAP_5699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19043__14 vssd1 vssd1 vccd1 vccd1 _19043__14/HI _19137_/A sky130_fd_sc_hd__conb_1
XFILLER_57_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16600_ _16659_/A vssd1 vssd1 vccd1 vccd1 _16600_/X sky130_fd_sc_hd__clkbuf_2
XTAP_4987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13812_ _12019_/B _13804_/X _13811_/X _12055_/B vssd1 vssd1 vccd1 vccd1 _13812_/X
+ sky130_fd_sc_hd__a22o_2
XFILLER_21_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17580_ _17580_/A vssd1 vssd1 vccd1 vccd1 _18957_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_217_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14792_ _18324_/Q _18288_/Q _14809_/S vssd1 vssd1 vccd1 vccd1 _14792_/X sky130_fd_sc_hd__mux2_1
XFILLER_63_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16531_ _18738_/Q _18702_/Q _16546_/S vssd1 vssd1 vccd1 vccd1 _16531_/X sky130_fd_sc_hd__mux2_1
XFILLER_16_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13743_ _13743_/A vssd1 vssd1 vccd1 vccd1 _13743_/X sky130_fd_sc_hd__buf_4
X_10955_ _09413_/A _09418_/D _10955_/S vssd1 vssd1 vccd1 vccd1 _10955_/X sky130_fd_sc_hd__mux2_1
XFILLER_216_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16462_ _18722_/Q _18686_/Q _16470_/S vssd1 vssd1 vccd1 vccd1 _16462_/X sky130_fd_sc_hd__mux2_1
XFILLER_32_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13674_ _18861_/Q _13522_/A _13586_/A _18864_/Q _13673_/X vssd1 vssd1 vccd1 vccd1
+ _13674_/X sky130_fd_sc_hd__a221o_1
X_10886_ _10757_/A _10881_/X _10885_/X _10616_/Y vssd1 vssd1 vccd1 vccd1 _10886_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_108_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18201_ _18908_/CLK _18201_/D vssd1 vssd1 vccd1 vccd1 _18201_/Q sky130_fd_sc_hd__dfxtp_1
X_15413_ _15442_/A _15417_/B vssd1 vssd1 vccd1 vccd1 _15413_/Y sky130_fd_sc_hd__nand2_1
XPHY_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_176_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12625_ _12627_/A vssd1 vssd1 vccd1 vccd1 _12653_/B sky130_fd_sc_hd__clkbuf_2
X_19181_ _19181_/A _09014_/Y vssd1 vssd1 vccd1 vccd1 io_out[19] sky130_fd_sc_hd__ebufn_8
XPHY_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_223_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16393_ _16392_/B _16391_/X _16392_/Y _16376_/X vssd1 vssd1 vccd1 vccd1 _18668_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_12_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_169_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18132_ _18972_/CLK _18132_/D vssd1 vssd1 vccd1 vccd1 _18132_/Q sky130_fd_sc_hd__dfxtp_1
X_15344_ _18456_/Q _18420_/Q _15356_/S vssd1 vssd1 vccd1 vccd1 _15344_/X sky130_fd_sc_hd__mux2_1
XFILLER_185_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12556_ _12556_/A _12556_/B vssd1 vssd1 vccd1 vccd1 _12557_/B sky130_fd_sc_hd__and2_1
XFILLER_156_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11507_ _11609_/A _11742_/A _11507_/C vssd1 vssd1 vccd1 vccd1 _11508_/B sky130_fd_sc_hd__or3_1
X_18063_ _18072_/CLK _18063_/D vssd1 vssd1 vccd1 vccd1 _18063_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_11_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15275_ _15303_/A _15275_/B vssd1 vssd1 vccd1 vccd1 _15275_/Y sky130_fd_sc_hd__nand2_1
X_12487_ _17909_/Q _12487_/B vssd1 vssd1 vccd1 vccd1 _12487_/Y sky130_fd_sc_hd__nor2_1
XFILLER_32_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17014_ _18852_/Q _18816_/Q _17026_/S vssd1 vssd1 vccd1 vccd1 _17014_/X sky130_fd_sc_hd__mux2_1
X_11438_ _11428_/B _11437_/X _11376_/A _11376_/B vssd1 vssd1 vccd1 vccd1 _11438_/X
+ sky130_fd_sc_hd__o211a_1
X_14226_ _14203_/X _14208_/X _14225_/Y vssd1 vssd1 vccd1 vccd1 _14226_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_67_1302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_217_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14157_ _18752_/Q _13568_/X _14155_/X _14156_/X vssd1 vssd1 vccd1 vccd1 _14157_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_193_1354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11369_ _11336_/A _11368_/Y _11297_/Y _11338_/A _11318_/A vssd1 vssd1 vccd1 vccd1
+ _11508_/C sky130_fd_sc_hd__o311ai_4
XFILLER_67_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_217_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13108_ _13108_/A vssd1 vssd1 vccd1 vccd1 _18014_/D sky130_fd_sc_hd__clkbuf_1
X_14088_ _14082_/X _14083_/X _14087_/X _11957_/B vssd1 vssd1 vccd1 vccd1 _14088_/X
+ sky130_fd_sc_hd__o31a_4
X_18965_ _18965_/CLK _18965_/D vssd1 vssd1 vccd1 vccd1 _18965_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_98_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_224_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_140_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17916_ _17919_/CLK _17916_/D vssd1 vssd1 vccd1 vccd1 _17916_/Q sky130_fd_sc_hd__dfxtp_1
X_13039_ _17992_/Q _13039_/B vssd1 vssd1 vccd1 vccd1 _13039_/X sky130_fd_sc_hd__or2_1
XFILLER_100_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18896_ _18899_/CLK _18896_/D vssd1 vssd1 vccd1 vccd1 _18896_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_224_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_227_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_230_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17847_ _17890_/CLK _17847_/D vssd1 vssd1 vccd1 vccd1 _17847_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_27_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17778_ _18191_/CLK _17778_/D vssd1 vssd1 vccd1 vccd1 _17778_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_214_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16729_ _18750_/Q _16732_/B _16728_/X _16724_/X vssd1 vssd1 vccd1 vccd1 _18750_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_62_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_223_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_1339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_228_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09201_ _18578_/Q _18577_/Q _18576_/Q vssd1 vssd1 vccd1 vccd1 _09203_/C sky130_fd_sc_hd__or3_4
Xclkbuf_leaf_56_wb_clk_i clkbuf_5_16_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18786_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_124_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09132_ _18821_/Q _18820_/Q _18819_/Q vssd1 vssd1 vccd1 vccd1 _09136_/A sky130_fd_sc_hd__or3_4
XFILLER_202_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09063_ _09072_/A _09069_/B _17825_/Q vssd1 vssd1 vccd1 vccd1 _09064_/A sky130_fd_sc_hd__and3_1
XFILLER_190_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_190_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_191_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09965_ _09965_/A vssd1 vssd1 vccd1 vccd1 _10338_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_131_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09896_ _10181_/A _09896_/B vssd1 vssd1 vccd1 vccd1 _09907_/B sky130_fd_sc_hd__or2_1
XTAP_4217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_217_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_3_3_0_wb_clk_i clkbuf_3_3_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_4_7_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_213_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10740_ _09993_/A _09153_/B _09148_/A _09143_/D _10858_/S _10764_/A vssd1 vssd1 vccd1
+ vccd1 _10740_/X sky130_fd_sc_hd__mux4_1
XFILLER_14_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_198_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_213_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10671_ _10753_/A _10671_/B _10671_/C vssd1 vssd1 vccd1 vccd1 _10671_/X sky130_fd_sc_hd__and3_1
XFILLER_199_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12410_ _12411_/B _17898_/Q vssd1 vssd1 vccd1 vccd1 _12412_/A sky130_fd_sc_hd__and2b_1
XFILLER_90_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_1294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13390_ _13346_/X _13389_/Y _13383_/A vssd1 vssd1 vccd1 vccd1 _18119_/D sky130_fd_sc_hd__a21boi_1
XFILLER_223_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12341_ _11479_/B _12347_/B _12340_/X _11822_/X vssd1 vssd1 vccd1 vccd1 _17886_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_142_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15060_ _18389_/Q _18353_/Q _15081_/S vssd1 vssd1 vccd1 vccd1 _15060_/X sky130_fd_sc_hd__mux2_1
XFILLER_5_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12272_ _12272_/A _12304_/A vssd1 vssd1 vccd1 vccd1 _12272_/X sky130_fd_sc_hd__and2_1
XFILLER_153_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14011_ _13846_/X _13867_/X _14010_/X _18167_/Q _14222_/A vssd1 vssd1 vccd1 vccd1
+ _14012_/B sky130_fd_sc_hd__o32a_2
XFILLER_49_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11223_ _11224_/A _11224_/C _11222_/Y vssd1 vssd1 vccd1 vccd1 _17817_/D sky130_fd_sc_hd__a21oi_1
XFILLER_49_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_122_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11154_ _15840_/A vssd1 vssd1 vccd1 vccd1 _12285_/A sky130_fd_sc_hd__buf_4
XFILLER_49_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10105_ _10017_/S _10102_/X _10104_/X _10076_/S vssd1 vssd1 vccd1 vccd1 _10105_/X
+ sky130_fd_sc_hd__a211o_1
X_18750_ _18752_/CLK _18750_/D vssd1 vssd1 vccd1 vccd1 _18750_/Q sky130_fd_sc_hd__dfxtp_2
X_15962_ _15962_/A _15993_/B vssd1 vssd1 vccd1 vccd1 _15971_/B sky130_fd_sc_hd__nor2_2
XFILLER_216_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11085_ _11951_/A vssd1 vssd1 vccd1 vccd1 _12023_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_110_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17701_ _14383_/B _13356_/B _14404_/X vssd1 vssd1 vccd1 vccd1 _17701_/Y sky130_fd_sc_hd__a21oi_1
XTAP_5463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14913_ _14935_/A _14913_/B vssd1 vssd1 vccd1 vccd1 _14913_/Y sky130_fd_sc_hd__nand2_1
X_10036_ _10036_/A vssd1 vssd1 vccd1 vccd1 _10036_/X sky130_fd_sc_hd__buf_4
X_18681_ _18683_/CLK _18681_/D vssd1 vssd1 vccd1 vccd1 _18681_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_5474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15893_ _18588_/Q _18552_/Q _15899_/S vssd1 vssd1 vccd1 vccd1 _15893_/X sky130_fd_sc_hd__mux2_1
XTAP_4740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17632_ _17571_/X _17623_/Y _17631_/X _17624_/Y _18971_/Q vssd1 vssd1 vccd1 vccd1
+ _17633_/B sky130_fd_sc_hd__a32o_1
XTAP_4773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14844_ _14849_/B _14842_/X _14843_/X _14839_/X vssd1 vssd1 vccd1 vccd1 _18300_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_224_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_189_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17563_ _17538_/A _17560_/Y _17561_/X _17562_/Y _18954_/Q vssd1 vssd1 vccd1 vccd1
+ _17564_/B sky130_fd_sc_hd__a32o_1
X_14775_ _14810_/A _14777_/B vssd1 vssd1 vccd1 vccd1 _14775_/Y sky130_fd_sc_hd__nand2_1
X_11987_ _11985_/B _11985_/D _11988_/C _12007_/A vssd1 vssd1 vccd1 vccd1 _12027_/C
+ sky130_fd_sc_hd__o211a_4
XFILLER_95_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_205_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16514_ _16578_/A vssd1 vssd1 vccd1 vccd1 _16652_/C sky130_fd_sc_hd__buf_2
XFILLER_16_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13726_ _18249_/Q _13723_/X _13725_/X _18231_/Q vssd1 vssd1 vccd1 vccd1 _13726_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_32_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17494_ _17501_/B _17492_/X _17493_/X _17478_/X vssd1 vssd1 vccd1 vccd1 _18936_/D
+ sky130_fd_sc_hd__o211a_1
X_10938_ _10443_/X _10918_/X _10924_/X _10270_/A _10937_/X vssd1 vssd1 vccd1 vccd1
+ _10938_/Y sky130_fd_sc_hd__a221oi_1
XFILLER_220_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19233_ _19233_/A _11018_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[33] sky130_fd_sc_hd__ebufn_8
X_16445_ _16450_/B _16442_/X _16444_/X _16437_/X vssd1 vssd1 vccd1 vccd1 _18681_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_189_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13657_ _13657_/A vssd1 vssd1 vccd1 vccd1 _13657_/X sky130_fd_sc_hd__buf_6
X_10869_ _09408_/A _09408_/B _09413_/C _09418_/B _10693_/X _10660_/X vssd1 vssd1 vccd1
+ vccd1 _10869_/X sky130_fd_sc_hd__mux4_1
XFILLER_32_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19164_ _19164_/A _09027_/Y vssd1 vssd1 vccd1 vccd1 io_out[2] sky130_fd_sc_hd__ebufn_8
X_12608_ _12608_/A vssd1 vssd1 vccd1 vccd1 _12637_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_223_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16376_ _16456_/A vssd1 vssd1 vccd1 vccd1 _16376_/X sky130_fd_sc_hd__clkbuf_2
XPHY_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13588_ _13588_/A vssd1 vssd1 vccd1 vccd1 _13588_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_185_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18115_ _19028_/CLK _18115_/D vssd1 vssd1 vccd1 vccd1 _18115_/Q sky130_fd_sc_hd__dfxtp_1
X_15327_ _16839_/A vssd1 vssd1 vccd1 vccd1 _15931_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_121_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12539_ _17918_/Q vssd1 vssd1 vccd1 vccd1 _12542_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_9_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_219_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18046_ _18052_/CLK _18046_/D vssd1 vssd1 vccd1 vccd1 _18046_/Q sky130_fd_sc_hd__dfxtp_1
X_15258_ _15263_/B _15256_/X _15257_/X _15244_/X vssd1 vssd1 vccd1 vccd1 _18402_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_32_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_172_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14209_ _18207_/Q _18206_/Q vssd1 vssd1 vccd1 vccd1 _14323_/C sky130_fd_sc_hd__or2_1
XFILLER_160_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15189_ _18421_/Q _18385_/Q _15198_/S vssd1 vssd1 vccd1 vccd1 _15189_/X sky130_fd_sc_hd__mux2_1
XFILLER_67_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_174_wb_clk_i clkbuf_5_11_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18993_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_63_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_103_wb_clk_i clkbuf_5_28_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18557_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_154_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_140_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09750_ _09749_/B _09749_/C _09802_/B vssd1 vssd1 vccd1 vccd1 _09751_/B sky130_fd_sc_hd__a21oi_1
X_18948_ _18950_/CLK _18948_/D vssd1 vssd1 vccd1 vccd1 _18948_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_113_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09681_ _10046_/A vssd1 vssd1 vccd1 vccd1 _09682_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_39_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18879_ _18907_/CLK _18879_/D vssd1 vssd1 vccd1 vccd1 _18879_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_66_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_215_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_214_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_120_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_1294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_223_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09115_ _18746_/Q _18745_/Q _18744_/Q vssd1 vssd1 vccd1 vccd1 _09119_/A sky130_fd_sc_hd__or3_4
XFILLER_13_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09046_ _09046_/A vssd1 vssd1 vccd1 vccd1 _09046_/Y sky130_fd_sc_hd__inv_2
XFILLER_136_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_1366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09948_ _09948_/A vssd1 vssd1 vccd1 vccd1 _14240_/B sky130_fd_sc_hd__buf_4
XTAP_4003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_20 _09214_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_31 _10600_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09879_ _09879_/A _09879_/B vssd1 vssd1 vccd1 vccd1 _09882_/A sky130_fd_sc_hd__xnor2_4
XTAP_4047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_42 _10940_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_213_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_53 _15840_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11910_ _11910_/A _11910_/B vssd1 vssd1 vccd1 vccd1 _11910_/Y sky130_fd_sc_hd__nor2_1
XTAP_3335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_64 _12510_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_75 _13576_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12890_ _17960_/Q _12890_/B vssd1 vssd1 vccd1 vccd1 _12895_/C sky130_fd_sc_hd__and2_1
XTAP_2601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_86 _13625_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XINSDIODE2_97 _13780_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11841_ _11513_/A _11840_/Y _11501_/X vssd1 vssd1 vccd1 vccd1 _11842_/C sky130_fd_sc_hd__o21ba_1
XTAP_2634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14560_ _17747_/A vssd1 vssd1 vccd1 vccd1 _14668_/A sky130_fd_sc_hd__buf_2
X_11772_ _11776_/B _11772_/B vssd1 vssd1 vccd1 vccd1 _11772_/X sky130_fd_sc_hd__or2_1
XFILLER_54_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_220_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_1304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_213_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_202_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10723_ _09148_/C _10737_/S _10722_/X _10743_/A vssd1 vssd1 vccd1 vccd1 _10723_/X
+ sky130_fd_sc_hd__o211a_1
X_13511_ _13667_/A vssd1 vssd1 vccd1 vccd1 _13734_/A sky130_fd_sc_hd__buf_6
XFILLER_18_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_207_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_144_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_202_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_1348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14491_ _18220_/Q _14491_/B vssd1 vssd1 vccd1 vccd1 _14492_/A sky130_fd_sc_hd__and2_1
XTAP_1988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16230_ _16252_/A vssd1 vssd1 vccd1 vccd1 _16230_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_220_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13442_ _13442_/A _13442_/B vssd1 vssd1 vccd1 vccd1 _13452_/B sky130_fd_sc_hd__xor2_1
XFILLER_16_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10654_ _10654_/A _12096_/B vssd1 vssd1 vccd1 vccd1 _10818_/B sky130_fd_sc_hd__nor2_4
XFILLER_174_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16161_ _16273_/A vssd1 vssd1 vccd1 vccd1 _16252_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_127_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13373_ _13346_/X _13372_/Y _13370_/B vssd1 vssd1 vccd1 vccd1 _18109_/D sky130_fd_sc_hd__a21boi_1
XFILLER_186_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10585_ _10962_/A _10582_/X _10584_/X _10086_/A vssd1 vssd1 vccd1 vccd1 _10585_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_155_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15112_ _15162_/A _15257_/B _15112_/C vssd1 vssd1 vccd1 vccd1 _15112_/X sky130_fd_sc_hd__or3_1
X_12324_ _11419_/X _12333_/C _12323_/X vssd1 vssd1 vccd1 vccd1 _12325_/B sky130_fd_sc_hd__a21oi_1
X_16092_ _16130_/A _16096_/B vssd1 vssd1 vccd1 vccd1 _16092_/Y sky130_fd_sc_hd__nand2_1
XFILLER_186_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_1_wb_clk_i clkbuf_5_0_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17926_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_5_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15043_ _15049_/B _15041_/X _15042_/X _15026_/X vssd1 vssd1 vccd1 vccd1 _18348_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_141_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12255_ _12270_/A vssd1 vssd1 vccd1 vccd1 _12276_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_170_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_190_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11206_ _11210_/A _11206_/B _11209_/B vssd1 vssd1 vccd1 vccd1 _11207_/A sky130_fd_sc_hd__and3_1
XFILLER_107_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12186_ _18989_/Q _18987_/Q _18105_/Q _18988_/Q vssd1 vssd1 vccd1 vccd1 _12401_/B
+ sky130_fd_sc_hd__or4_4
XFILLER_69_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18802_ _18806_/CLK _18802_/D vssd1 vssd1 vccd1 vccd1 _18802_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_123_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11137_ _11253_/A _11196_/B _11149_/S vssd1 vssd1 vccd1 vccd1 _11138_/A sky130_fd_sc_hd__mux2_1
XFILLER_228_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16994_ _18847_/Q _18811_/Q _17005_/S vssd1 vssd1 vccd1 vccd1 _16994_/X sky130_fd_sc_hd__mux2_1
XFILLER_95_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18733_ _18765_/CLK _18733_/D vssd1 vssd1 vccd1 vccd1 _18733_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_27_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15945_ _18600_/Q _18564_/Q _15963_/S vssd1 vssd1 vccd1 vccd1 _15945_/X sky130_fd_sc_hd__mux2_1
XTAP_5260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11068_ _11334_/B vssd1 vssd1 vccd1 vccd1 _11368_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_62_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_225_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10019_ _09114_/B _09109_/B _10019_/S vssd1 vssd1 vccd1 vccd1 _10019_/X sky130_fd_sc_hd__mux2_1
XFILLER_23_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18664_ _18696_/CLK _18664_/D vssd1 vssd1 vccd1 vccd1 _18664_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_114_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15876_ _15876_/A _15876_/B vssd1 vssd1 vccd1 vccd1 _15876_/Y sky130_fd_sc_hd__nand2_1
XTAP_4570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_221_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_1264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17615_ _17615_/A vssd1 vssd1 vccd1 vccd1 _18965_/D sky130_fd_sc_hd__clkbuf_1
X_14827_ _14875_/A _14827_/B vssd1 vssd1 vccd1 vccd1 _14827_/Y sky130_fd_sc_hd__nand2_1
XFILLER_64_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18595_ _18608_/CLK _18595_/D vssd1 vssd1 vccd1 vccd1 _18595_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_184_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17546_ _17549_/A _17549_/B vssd1 vssd1 vccd1 vccd1 _17547_/A sky130_fd_sc_hd__or2_1
X_14758_ _14778_/A vssd1 vssd1 vccd1 vccd1 _14758_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_32_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13709_ _18741_/Q _13546_/A _13701_/X _13708_/X vssd1 vssd1 vccd1 vccd1 _13709_/X
+ sky130_fd_sc_hd__a211o_1
X_17477_ _17512_/A _17477_/B vssd1 vssd1 vccd1 vccd1 _17477_/Y sky130_fd_sc_hd__nand2_1
X_14689_ _16962_/A vssd1 vssd1 vccd1 vccd1 _15279_/B sky130_fd_sc_hd__buf_6
XFILLER_225_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19216_ _19216_/A _08969_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[16] sky130_fd_sc_hd__ebufn_8
X_16428_ _18713_/Q _18677_/Q _16449_/S vssd1 vssd1 vccd1 vccd1 _16428_/X sky130_fd_sc_hd__mux2_1
XFILLER_177_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19147_ _19147_/A _09043_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[17] sky130_fd_sc_hd__ebufn_8
XFILLER_9_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16359_ _16364_/B _16357_/X _16358_/X _16354_/X vssd1 vssd1 vccd1 vccd1 _18660_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_117_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18029_ _18087_/CLK _18029_/D vssd1 vssd1 vccd1 vccd1 _18029_/Q sky130_fd_sc_hd__dfxtp_1
X_19079__50 vssd1 vssd1 vccd1 vccd1 _19079__50/HI _19187_/A sky130_fd_sc_hd__conb_1
XFILLER_132_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09802_ _17982_/Q _09802_/B vssd1 vssd1 vccd1 vccd1 _09806_/A sky130_fd_sc_hd__xnor2_1
XFILLER_86_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_1260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09733_ _18102_/Q vssd1 vssd1 vccd1 vccd1 _09743_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_41_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09664_ _09664_/A _09664_/B vssd1 vssd1 vccd1 vccd1 _12072_/B sky130_fd_sc_hd__xnor2_2
XFILLER_131_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_216_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09595_ _09723_/A _09722_/B _09594_/X vssd1 vssd1 vccd1 vccd1 _09726_/A sky130_fd_sc_hd__a21o_2
Xclkbuf_leaf_71_wb_clk_i clkbuf_5_20_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18663_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_1207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_211_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_190 _09109_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_1280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_210_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10370_ _10368_/X _10369_/X _10370_/S vssd1 vssd1 vccd1 vccd1 _10370_/X sky130_fd_sc_hd__mux2_1
XFILLER_100_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_136_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09029_ _09029_/A vssd1 vssd1 vccd1 vccd1 _09034_/A sky130_fd_sc_hd__buf_12
XFILLER_191_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12040_ _12120_/A _11920_/B _12035_/X _12039_/X vssd1 vssd1 vccd1 vccd1 _12040_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_123_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_5_24_0_wb_clk_i clkbuf_5_25_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_5_24_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_172_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_219_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_1333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13991_ _18382_/Q _13651_/X _13985_/X _13990_/X vssd1 vssd1 vccd1 vccd1 _13991_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_213_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_1366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15730_ _15754_/A _15730_/B vssd1 vssd1 vccd1 vccd1 _15730_/Y sky130_fd_sc_hd__nand2_1
XFILLER_58_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_219_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_218_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12942_ _17972_/Q vssd1 vssd1 vccd1 vccd1 _13368_/A sky130_fd_sc_hd__buf_2
XFILLER_58_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15661_ _15694_/A _15661_/B vssd1 vssd1 vccd1 vccd1 _15661_/Y sky130_fd_sc_hd__nand2_1
XTAP_2420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12873_ _12877_/C _12873_/B vssd1 vssd1 vccd1 vccd1 _17954_/D sky130_fd_sc_hd__nor2_1
XFILLER_74_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17400_ _17400_/A vssd1 vssd1 vccd1 vccd1 _17400_/X sky130_fd_sc_hd__clkbuf_2
XTAP_3187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14612_ _14612_/A vssd1 vssd1 vccd1 vccd1 _14612_/X sky130_fd_sc_hd__buf_2
XTAP_3198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18380_ _18380_/CLK _18380_/D vssd1 vssd1 vccd1 vccd1 _18380_/Q sky130_fd_sc_hd__dfxtp_2
X_11824_ _11824_/A vssd1 vssd1 vccd1 vccd1 _11826_/A sky130_fd_sc_hd__inv_2
XTAP_2464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15592_ _15594_/B _15590_/X _15591_/Y _15575_/X vssd1 vssd1 vccd1 vccd1 _18478_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_1730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17331_ _17331_/A vssd1 vssd1 vccd1 vccd1 _17376_/C sky130_fd_sc_hd__clkbuf_1
X_14543_ _15649_/A vssd1 vssd1 vccd1 vccd1 _17544_/A sky130_fd_sc_hd__buf_2
XTAP_1763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11755_ _11727_/A _11737_/B _11767_/A vssd1 vssd1 vccd1 vccd1 _11756_/S sky130_fd_sc_hd__o21ai_1
XTAP_1774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_222_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10706_ _13000_/A _10706_/B vssd1 vssd1 vccd1 vccd1 _10843_/B sky130_fd_sc_hd__xnor2_4
XFILLER_81_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17262_ _18914_/Q _18878_/Q _17262_/S vssd1 vssd1 vccd1 vccd1 _17262_/X sky130_fd_sc_hd__mux2_1
XFILLER_140_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14474_ _18212_/Q _14480_/B vssd1 vssd1 vccd1 vccd1 _14475_/A sky130_fd_sc_hd__and2_1
XFILLER_105_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11686_ _17851_/Q vssd1 vssd1 vccd1 vccd1 _11703_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_144_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19001_ _19026_/CLK _19001_/D vssd1 vssd1 vccd1 vccd1 _19001_/Q sky130_fd_sc_hd__dfxtp_1
X_16213_ _16265_/A _16217_/B vssd1 vssd1 vccd1 vccd1 _16213_/Y sky130_fd_sc_hd__nand2_1
XFILLER_179_1208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13425_ _12055_/C _13710_/C _13435_/B vssd1 vssd1 vccd1 vccd1 _13426_/B sky130_fd_sc_hd__o21ai_4
XFILLER_220_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10637_ _10654_/A _12096_/B vssd1 vssd1 vccd1 vccd1 _10667_/A sky130_fd_sc_hd__or2_1
X_17193_ _17193_/A _17483_/B _17234_/C vssd1 vssd1 vccd1 vccd1 _17193_/X sky130_fd_sc_hd__or3_1
XFILLER_31_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16144_ _16147_/B _16141_/X _16143_/Y _16139_/X vssd1 vssd1 vccd1 vccd1 _18610_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_155_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10568_ _10568_/A vssd1 vssd1 vccd1 vccd1 _10568_/X sky130_fd_sc_hd__buf_2
X_13356_ _17704_/A _13356_/B vssd1 vssd1 vccd1 vccd1 _13356_/Y sky130_fd_sc_hd__nor2_1
XFILLER_170_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_154_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12307_ _11339_/D _12292_/B _11323_/A vssd1 vssd1 vccd1 vccd1 _12307_/Y sky130_fd_sc_hd__a21oi_1
X_16075_ _16082_/B _16071_/X _16073_/X _16074_/X vssd1 vssd1 vccd1 vccd1 _18594_/D
+ sky130_fd_sc_hd__o211a_1
X_13287_ _18013_/Q _18012_/Q _18015_/Q _18014_/Q vssd1 vssd1 vccd1 vccd1 _13291_/A
+ sky130_fd_sc_hd__or4_1
XFILLER_5_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10499_ _10932_/A _10496_/Y _10498_/X _12031_/A _10456_/A vssd1 vssd1 vccd1 vccd1
+ _10499_/X sky130_fd_sc_hd__a311o_1
XFILLER_216_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15026_ _15083_/A vssd1 vssd1 vccd1 vccd1 _15026_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_155_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12238_ _11603_/A _12235_/Y _12258_/C _12219_/X vssd1 vssd1 vccd1 vccd1 _17858_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_107_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12169_ _12169_/A _12169_/B vssd1 vssd1 vccd1 vccd1 _12180_/A sky130_fd_sc_hd__nor2_1
XFILLER_9_1349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_116_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16977_ _17012_/A vssd1 vssd1 vccd1 vccd1 _17107_/B sky130_fd_sc_hd__buf_2
XFILLER_96_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_231_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput5 io_in[27] vssd1 vssd1 vccd1 vccd1 input5/X sky130_fd_sc_hd__clkbuf_2
XFILLER_65_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15928_ _15942_/A _15928_/B vssd1 vssd1 vccd1 vccd1 _15928_/Y sky130_fd_sc_hd__nand2_1
X_18716_ _18752_/CLK _18716_/D vssd1 vssd1 vccd1 vccd1 _18716_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_5090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18647_ _18683_/CLK _18647_/D vssd1 vssd1 vccd1 vccd1 _18647_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_65_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15859_ _18580_/Q _18544_/Q _15859_/S vssd1 vssd1 vccd1 vccd1 _15859_/X sky130_fd_sc_hd__mux2_1
XFILLER_188_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_224_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09380_ _18401_/Q _18400_/Q _18399_/Q vssd1 vssd1 vccd1 vccd1 _09381_/D sky130_fd_sc_hd__or3_4
XFILLER_24_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18578_ _18593_/CLK _18578_/D vssd1 vssd1 vccd1 vccd1 _18578_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_51_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_212_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_224_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17529_ _17534_/B _17527_/X _17528_/X _17517_/X vssd1 vssd1 vccd1 vccd1 _18945_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_33_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_221_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_195_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_142_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_1208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09716_ _10085_/S vssd1 vssd1 vccd1 vccd1 _10065_/A sky130_fd_sc_hd__buf_6
XFILLER_132_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_228_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_215_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09647_ _09647_/A _09647_/B vssd1 vssd1 vccd1 vccd1 _09684_/B sky130_fd_sc_hd__xnor2_1
XFILLER_216_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09578_ _09580_/A _09578_/B vssd1 vssd1 vccd1 vccd1 _09600_/B sky130_fd_sc_hd__xnor2_1
XTAP_1037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11540_ _11735_/A _11593_/A _11770_/C _11654_/B vssd1 vssd1 vccd1 vccd1 _11546_/A
+ sky130_fd_sc_hd__or4b_1
XFILLER_51_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_168_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_206_wb_clk_i clkbuf_5_6_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18965_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_183_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11471_ _17886_/Q vssd1 vssd1 vccd1 vccd1 _11472_/A sky130_fd_sc_hd__inv_2
XFILLER_52_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13210_ _13210_/A vssd1 vssd1 vccd1 vccd1 _13467_/A sky130_fd_sc_hd__buf_6
X_10422_ _10422_/A vssd1 vssd1 vccd1 vccd1 _14307_/A sky130_fd_sc_hd__buf_2
X_14190_ _18210_/Q vssd1 vssd1 vccd1 vccd1 _14470_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_178_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10353_ _12128_/A _10347_/X _10352_/X _09921_/X vssd1 vssd1 vccd1 vccd1 _10353_/X
+ sky130_fd_sc_hd__o211a_1
X_13141_ _13141_/A vssd1 vssd1 vccd1 vccd1 _18029_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_87_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13072_ _18152_/Q _13269_/B vssd1 vssd1 vccd1 vccd1 _13072_/X sky130_fd_sc_hd__or2_1
XFILLER_151_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10284_ _09930_/X _10282_/X _10283_/X _10278_/X vssd1 vssd1 vccd1 vccd1 _10288_/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_152_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16900_ _18827_/Q _18791_/Q _16900_/S vssd1 vssd1 vccd1 vccd1 _16900_/X sky130_fd_sc_hd__mux2_1
XFILLER_2_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12023_ _12023_/A _12023_/B vssd1 vssd1 vccd1 vccd1 _12023_/Y sky130_fd_sc_hd__nor2_1
X_17880_ _17883_/CLK _17880_/D vssd1 vssd1 vccd1 vccd1 _17880_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_215_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16831_ _18812_/Q _18776_/Q _16842_/S vssd1 vssd1 vccd1 vccd1 _16831_/X sky130_fd_sc_hd__mux2_1
XFILLER_76_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16762_ _18796_/Q _18760_/Q _16762_/S vssd1 vssd1 vccd1 vccd1 _16762_/X sky130_fd_sc_hd__mux2_1
X_13974_ _18286_/Q _13742_/X _13766_/X _18268_/Q vssd1 vssd1 vccd1 vccd1 _13974_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_4_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18501_ _18532_/CLK _18501_/D vssd1 vssd1 vccd1 vccd1 _18501_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_150_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15713_ _15719_/B _15711_/X _15712_/X _15700_/X vssd1 vssd1 vccd1 vccd1 _18507_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_185_1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12925_ _18153_/Q _12925_/B vssd1 vssd1 vccd1 vccd1 _12927_/A sky130_fd_sc_hd__or2_1
X_16693_ _16699_/B _16690_/X _16692_/X _16683_/X vssd1 vssd1 vccd1 vccd1 _18741_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_47_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18432_ _18432_/CLK _18432_/D vssd1 vssd1 vccd1 vccd1 _18432_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_185_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15644_ _15885_/A vssd1 vssd1 vccd1 vccd1 _15691_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_18_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12856_ _12816_/X _12857_/C _12855_/Y vssd1 vssd1 vccd1 vccd1 _17949_/D sky130_fd_sc_hd__a21oi_1
XTAP_2261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18363_ _18367_/CLK _18363_/D vssd1 vssd1 vccd1 vccd1 _18363_/Q sky130_fd_sc_hd__dfxtp_2
X_11807_ _11807_/A _11937_/C vssd1 vssd1 vccd1 vccd1 _11807_/X sky130_fd_sc_hd__or2_1
XTAP_2294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15575_ _15616_/A vssd1 vssd1 vccd1 vccd1 _15575_/X sky130_fd_sc_hd__clkbuf_2
XTAP_1560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12787_ _13082_/A _13066_/C _12786_/X _12318_/X vssd1 vssd1 vccd1 vccd1 _17943_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_203_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17314_ _17336_/A _17314_/B vssd1 vssd1 vccd1 vccd1 _17314_/Y sky130_fd_sc_hd__nand2_1
XFILLER_187_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14526_ _14704_/C _14526_/B vssd1 vssd1 vccd1 vccd1 _14598_/A sky130_fd_sc_hd__or2_4
XFILLER_186_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18294_ _18296_/CLK _18294_/D vssd1 vssd1 vccd1 vccd1 _18294_/Q sky130_fd_sc_hd__dfxtp_1
X_11738_ _17914_/Q _11737_/B _17913_/Q vssd1 vssd1 vccd1 vccd1 _11747_/A sky130_fd_sc_hd__o21ai_2
XFILLER_226_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_230_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17245_ _17256_/A _17528_/B _17256_/C vssd1 vssd1 vccd1 vccd1 _17245_/X sky130_fd_sc_hd__or3_1
XFILLER_35_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14457_ _18205_/Q _14457_/B _14457_/C vssd1 vssd1 vccd1 vccd1 _14458_/A sky130_fd_sc_hd__and3_1
X_11669_ _11669_/A _11669_/B _11669_/C vssd1 vssd1 vccd1 vccd1 _11669_/X sky130_fd_sc_hd__or3_1
X_13408_ _18130_/Q _11021_/X _13337_/X _13395_/X vssd1 vssd1 vccd1 vccd1 _18130_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_162_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17176_ _18892_/Q _18856_/Q _17199_/S vssd1 vssd1 vccd1 vccd1 _17176_/X sky130_fd_sc_hd__mux2_1
X_14388_ _18189_/Q _14386_/Y _14387_/X vssd1 vssd1 vccd1 vccd1 _18189_/D sky130_fd_sc_hd__o21ba_1
XFILLER_196_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16127_ _16127_/A vssd1 vssd1 vccd1 vccd1 _16181_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_192_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13339_ _17768_/B vssd1 vssd1 vccd1 vccd1 _13339_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_51_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_227_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16058_ _16127_/A vssd1 vssd1 vccd1 vccd1 _16205_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_157_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19049__20 vssd1 vssd1 vccd1 vccd1 _19049__20/HI _19143_/A sky130_fd_sc_hd__conb_1
XFILLER_97_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15009_ _18340_/Q _15012_/B _15008_/Y _15004_/X vssd1 vssd1 vccd1 vccd1 _18340_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_116_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_123_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_229_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09501_ _18199_/Q _09501_/B vssd1 vssd1 vccd1 vccd1 _09502_/B sky130_fd_sc_hd__or2_1
XFILLER_53_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09432_ _09470_/A _09432_/B _09432_/C vssd1 vssd1 vccd1 vccd1 _09435_/B sky130_fd_sc_hd__and3b_1
XFILLER_164_1307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_227_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_198_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09363_ _18302_/Q _18301_/Q _18300_/Q vssd1 vssd1 vccd1 vccd1 _09365_/C sky130_fd_sc_hd__or3_2
XFILLER_12_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_212_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09294_ _09294_/A _09294_/B _09294_/C _09294_/D vssd1 vssd1 vccd1 vccd1 _09294_/X
+ sky130_fd_sc_hd__and4_1
XFILLER_123_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_221_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_197_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_193_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_173_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_1207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10971_ _18230_/Q _18229_/Q _14515_/B vssd1 vssd1 vccd1 vccd1 _13417_/B sky130_fd_sc_hd__nor3_2
XFILLER_46_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12710_ _17938_/Q _12707_/X _11218_/X vssd1 vssd1 vccd1 vccd1 _12710_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_189_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_216_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13690_ _18609_/Q _13594_/A _13535_/A _18591_/Q vssd1 vssd1 vccd1 vccd1 _13690_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_188_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_203_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12641_ _12640_/A _12640_/B _12591_/X vssd1 vssd1 vccd1 vccd1 _12641_/X sky130_fd_sc_hd__o21a_1
XFILLER_70_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_231_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15360_ _15415_/A vssd1 vssd1 vccd1 vccd1 _15388_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_196_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_168_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12572_ _17924_/Q _12574_/B vssd1 vssd1 vccd1 vccd1 _12573_/A sky130_fd_sc_hd__nand2_1
XFILLER_180_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14311_ _14311_/A _14311_/B vssd1 vssd1 vccd1 vccd1 _14321_/A sky130_fd_sc_hd__and2_1
XFILLER_184_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11523_ _11390_/A _11515_/Y _11522_/X _11525_/B vssd1 vssd1 vccd1 vccd1 _11523_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_11_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15291_ _15370_/A vssd1 vssd1 vccd1 vccd1 _15451_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_183_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_1268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17030_ _17078_/A vssd1 vssd1 vccd1 vccd1 _17055_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_8_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14242_ _14219_/X _14234_/Y _14241_/X _14222_/Y vssd1 vssd1 vccd1 vccd1 _14242_/X
+ sky130_fd_sc_hd__a211o_1
X_11454_ _11546_/B _11482_/A vssd1 vssd1 vccd1 vccd1 _11455_/D sky130_fd_sc_hd__and2_1
XFILLER_137_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10405_ _09930_/X _10372_/X _10395_/X _10366_/X _10404_/Y vssd1 vssd1 vccd1 vccd1
+ _10405_/X sky130_fd_sc_hd__a221o_1
XFILLER_194_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14173_ _18599_/Q _13546_/X _14169_/X _14172_/X vssd1 vssd1 vccd1 vccd1 _14173_/X
+ sky130_fd_sc_hd__a211o_1
X_11385_ _11385_/A _11385_/B vssd1 vssd1 vccd1 vccd1 _11385_/X sky130_fd_sc_hd__and2_1
XFILLER_152_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13124_ _13124_/A vssd1 vssd1 vccd1 vccd1 _18021_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_194_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10336_ _10328_/X _10335_/X _09983_/B vssd1 vssd1 vccd1 vccd1 _10336_/X sky130_fd_sc_hd__o21a_1
XFILLER_98_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18981_ _18986_/CLK _18981_/D vssd1 vssd1 vccd1 vccd1 _18981_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_140_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_152_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10267_ _09370_/A _09360_/B _09360_/A _09365_/C _10231_/X _10236_/X vssd1 vssd1 vccd1
+ vccd1 _10267_/X sky130_fd_sc_hd__mux4_2
XFILLER_3_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13055_ _13080_/A _13055_/B vssd1 vssd1 vccd1 vccd1 _13055_/X sky130_fd_sc_hd__or2_1
X_17932_ _17933_/CLK _17932_/D vssd1 vssd1 vccd1 vccd1 _17932_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_87_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12006_ _12006_/A _12006_/B _12018_/A vssd1 vssd1 vccd1 vccd1 _12048_/A sky130_fd_sc_hd__and3_1
X_17863_ _19032_/CLK _17863_/D vssd1 vssd1 vccd1 vccd1 _17863_/Q sky130_fd_sc_hd__dfxtp_1
X_10198_ _10215_/A _10201_/B vssd1 vssd1 vccd1 vccd1 _10202_/A sky130_fd_sc_hd__nor2_1
XFILLER_38_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_226_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16814_ _18772_/Q _16815_/B _16813_/Y _16800_/X vssd1 vssd1 vccd1 vccd1 _18772_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_19_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17794_ _17824_/CLK _17794_/D vssd1 vssd1 vccd1 vccd1 _17794_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_93_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16745_ _16745_/A _16745_/B vssd1 vssd1 vccd1 vccd1 _16755_/B sky130_fd_sc_hd__nor2_1
X_13957_ _18649_/Q _13560_/A _13654_/X _18640_/Q _13956_/X vssd1 vssd1 vccd1 vccd1
+ _13957_/X sky130_fd_sc_hd__a221o_1
XFILLER_35_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_199_wb_clk_i _18176_/CLK vssd1 vssd1 vccd1 vccd1 _18182_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_62_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12908_ _17966_/Q _12908_/B vssd1 vssd1 vccd1 vccd1 _12913_/C sky130_fd_sc_hd__and2_1
X_16676_ _16766_/A vssd1 vssd1 vccd1 vccd1 _16694_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_61_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13888_ _18982_/Q _13657_/X _13886_/X _13887_/X vssd1 vssd1 vccd1 vccd1 _13888_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_207_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_128_wb_clk_i clkbuf_5_24_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18393_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_18415_ _18416_/CLK _18415_/D vssd1 vssd1 vccd1 vccd1 _18415_/Q sky130_fd_sc_hd__dfxtp_2
X_15627_ _15678_/A _15921_/B _15666_/C vssd1 vssd1 vccd1 vccd1 _15627_/X sky130_fd_sc_hd__or3_1
XFILLER_146_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_222_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12839_ _12839_/A _12888_/B vssd1 vssd1 vccd1 vccd1 _12840_/A sky130_fd_sc_hd__and2_1
XTAP_2080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_222_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18346_ _18346_/CLK _18346_/D vssd1 vssd1 vccd1 vccd1 _18346_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_61_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15558_ _15570_/A _15558_/B vssd1 vssd1 vccd1 vccd1 _15558_/Y sky130_fd_sc_hd__nand2_1
XTAP_1390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_187_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14509_ _14507_/A _14355_/B _14515_/C vssd1 vssd1 vccd1 vccd1 _14510_/C sky130_fd_sc_hd__a21bo_1
X_18277_ _18278_/CLK _18277_/D vssd1 vssd1 vccd1 vccd1 _18277_/Q sky130_fd_sc_hd__dfxtp_1
X_15489_ _15529_/A vssd1 vssd1 vccd1 vccd1 _15548_/B sky130_fd_sc_hd__buf_2
XFILLER_175_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17228_ _17228_/A vssd1 vssd1 vccd1 vccd1 _17468_/A sky130_fd_sc_hd__buf_2
XFILLER_147_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17159_ _18888_/Q _18852_/Q _17172_/S vssd1 vssd1 vccd1 vccd1 _17159_/X sky130_fd_sc_hd__mux2_1
Xclkbuf_4_5_0_wb_clk_i clkbuf_4_5_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_4_5_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_196_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09981_ _09981_/A vssd1 vssd1 vccd1 vccd1 _09981_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_107_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08932_ _08935_/A vssd1 vssd1 vccd1 vccd1 _08932_/Y sky130_fd_sc_hd__inv_2
XFILLER_170_1311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_168_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_225_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09415_ _18326_/Q _18325_/Q _18324_/Q vssd1 vssd1 vccd1 vccd1 _09418_/B sky130_fd_sc_hd__or3_2
XFILLER_52_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_209_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_197_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09346_ _18431_/Q _18430_/Q _18429_/Q vssd1 vssd1 vccd1 vccd1 _09349_/B sky130_fd_sc_hd__or3_4
XFILLER_12_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09277_ _09277_/A _09277_/B _09277_/C _09277_/D vssd1 vssd1 vccd1 vccd1 _09288_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_166_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11170_ _12361_/A vssd1 vssd1 vccd1 vccd1 _17661_/A sky130_fd_sc_hd__buf_6
XFILLER_162_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10121_ _10133_/A _10121_/B vssd1 vssd1 vccd1 vccd1 _10131_/A sky130_fd_sc_hd__or2_2
XFILLER_121_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_216_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10052_ _10069_/A _10050_/X _10051_/X _10086_/A _10029_/S vssd1 vssd1 vccd1 vccd1
+ _10053_/B sky130_fd_sc_hd__a221o_1
XTAP_5634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_216_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14860_ _18304_/Q _14861_/B _14858_/Y _14859_/X vssd1 vssd1 vccd1 vccd1 _18304_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_5689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13811_ _18408_/Q _13759_/A _13780_/A _18399_/Q _13810_/X vssd1 vssd1 vccd1 vccd1
+ _13811_/X sky130_fd_sc_hd__a221o_1
XFILLER_21_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14791_ _14812_/A vssd1 vssd1 vccd1 vccd1 _14809_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_95_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_217_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16530_ _16621_/A vssd1 vssd1 vccd1 vccd1 _16546_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_21_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_216_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13742_ _13785_/A vssd1 vssd1 vccd1 vccd1 _13742_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_17_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10954_ _09418_/A _09413_/D _09408_/D _09418_/C _09683_/X _09709_/X vssd1 vssd1 vccd1
+ vccd1 _10954_/X sky130_fd_sc_hd__mux4_1
XFILLER_43_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_221_wb_clk_i _17803_/CLK vssd1 vssd1 vccd1 vccd1 _17851_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_231_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16461_ _16464_/B _16458_/X _16460_/Y _16456_/X vssd1 vssd1 vccd1 vccd1 _18685_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_44_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13673_ _18858_/Q _13666_/X _13669_/X _13672_/X vssd1 vssd1 vccd1 vccd1 _13673_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_95_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10885_ _10648_/X _10882_/X _10884_/X _10700_/S vssd1 vssd1 vccd1 vccd1 _10885_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_43_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18200_ _18203_/CLK _18200_/D vssd1 vssd1 vccd1 vccd1 _18200_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_231_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_223_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15412_ _18472_/Q _18436_/Q _15412_/S vssd1 vssd1 vccd1 vccd1 _15412_/X sky130_fd_sc_hd__mux2_1
XPHY_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19180_ _19180_/A _09013_/Y vssd1 vssd1 vccd1 vccd1 io_out[18] sky130_fd_sc_hd__ebufn_8
X_12624_ _17930_/Q vssd1 vssd1 vccd1 vccd1 _12627_/A sky130_fd_sc_hd__inv_2
XPHY_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16392_ _16392_/A _16392_/B vssd1 vssd1 vccd1 vccd1 _16392_/Y sky130_fd_sc_hd__nand2_1
XPHY_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_223_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18131_ _18972_/CLK _18131_/D vssd1 vssd1 vccd1 vccd1 _18131_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_106_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15343_ _15944_/A _15393_/B vssd1 vssd1 vccd1 vccd1 _15352_/B sky130_fd_sc_hd__nor2_1
XFILLER_196_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12555_ _12574_/B _17918_/Q _12535_/A _12535_/B _12543_/X vssd1 vssd1 vccd1 vccd1
+ _12556_/B sky130_fd_sc_hd__a221o_1
XFILLER_11_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_223_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18062_ _18072_/CLK _18062_/D vssd1 vssd1 vccd1 vccd1 _18062_/Q sky130_fd_sc_hd__dfxtp_1
X_11506_ _11654_/C _11506_/B _11497_/B vssd1 vssd1 vccd1 vccd1 _11507_/C sky130_fd_sc_hd__or3b_1
X_15274_ _18443_/Q _18407_/Q _15285_/S vssd1 vssd1 vccd1 vccd1 _15274_/X sky130_fd_sc_hd__mux2_1
X_12486_ _17909_/Q _12486_/B vssd1 vssd1 vccd1 vccd1 _12492_/A sky130_fd_sc_hd__and2_1
XFILLER_138_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17013_ _17446_/A _17070_/B vssd1 vssd1 vccd1 vccd1 _17023_/B sky130_fd_sc_hd__nor2_2
XFILLER_32_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14225_ _14219_/X _14222_/Y _14224_/Y vssd1 vssd1 vccd1 vccd1 _14225_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_208_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11437_ _11423_/A _12316_/B _11431_/Y vssd1 vssd1 vccd1 vccd1 _11437_/X sky130_fd_sc_hd__o21a_1
XFILLER_67_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_125_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14156_ _18767_/Q _13940_/X _14030_/X _18764_/Q vssd1 vssd1 vccd1 vccd1 _14156_/X
+ sky130_fd_sc_hd__a22o_1
X_11368_ _11368_/A _11368_/B vssd1 vssd1 vccd1 vccd1 _11368_/Y sky130_fd_sc_hd__nand2_1
XFILLER_28_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_193_1366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13107_ _13107_/A _18015_/Q vssd1 vssd1 vccd1 vccd1 _13108_/A sky130_fd_sc_hd__and2_1
X_10319_ _09969_/X _10316_/X _10318_/X _10356_/A vssd1 vssd1 vccd1 vccd1 _10319_/X
+ sky130_fd_sc_hd__a211o_1
X_14087_ _18464_/Q _13834_/X _14085_/X _14086_/X vssd1 vssd1 vccd1 vccd1 _14087_/X
+ sky130_fd_sc_hd__a211o_1
X_18964_ _18970_/CLK _18964_/D vssd1 vssd1 vccd1 vccd1 _18964_/Q sky130_fd_sc_hd__dfxtp_2
X_11299_ _11337_/A _12023_/B _11296_/Y _11297_/Y _11298_/X vssd1 vssd1 vccd1 vccd1
+ _11301_/A sky130_fd_sc_hd__a32o_1
XFILLER_79_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_224_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_230_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13038_ _13005_/A _13025_/X _13036_/X _13037_/X vssd1 vssd1 vccd1 vccd1 _17991_/D
+ sky130_fd_sc_hd__o211a_1
X_17915_ _18960_/CLK _17915_/D vssd1 vssd1 vccd1 vccd1 _17915_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_140_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18895_ _18899_/CLK _18895_/D vssd1 vssd1 vccd1 vccd1 _18895_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_94_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17846_ _18163_/CLK _17846_/D vssd1 vssd1 vccd1 vccd1 _17846_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_14_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14989_ _15042_/A _15279_/B _14989_/C vssd1 vssd1 vccd1 vccd1 _14989_/X sky130_fd_sc_hd__or3_1
X_17777_ _19035_/Q _12246_/Y _12178_/X vssd1 vssd1 vccd1 vccd1 _19035_/D sky130_fd_sc_hd__o21a_1
XFILLER_81_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16728_ _16736_/A _16880_/B _16773_/C vssd1 vssd1 vccd1 vccd1 _16728_/X sky130_fd_sc_hd__or3_1
XFILLER_35_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_222_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_223_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16659_ _16659_/A vssd1 vssd1 vccd1 vccd1 _16659_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_50_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19036__7 vssd1 vssd1 vccd1 vccd1 _19036__7/HI _19130_/A sky130_fd_sc_hd__conb_1
XFILLER_222_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09200_ _18563_/Q _18562_/Q _18561_/Q vssd1 vssd1 vccd1 vccd1 _09203_/B sky130_fd_sc_hd__or3_4
XFILLER_50_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_176_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09131_ _09131_/A _09131_/B _09131_/C _09131_/D vssd1 vssd1 vccd1 vccd1 _09137_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_124_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18329_ _18346_/CLK _18329_/D vssd1 vssd1 vccd1 vccd1 _18329_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_147_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_198_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09062_ _17837_/Q vssd1 vssd1 vccd1 vccd1 _09069_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_135_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_25_wb_clk_i clkbuf_5_6_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18926_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_150_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_144_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09964_ _10388_/A _09964_/B vssd1 vssd1 vccd1 vccd1 _09964_/X sky130_fd_sc_hd__or2_1
XFILLER_134_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09895_ _09965_/A vssd1 vssd1 vccd1 vccd1 _09895_/X sky130_fd_sc_hd__clkbuf_4
XTAP_960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_225_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_230_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_198_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10670_ _09344_/B _09354_/C _10391_/A _10389_/A _10811_/A _10882_/S vssd1 vssd1 vccd1
+ vccd1 _10671_/C sky130_fd_sc_hd__mux4_1
XFILLER_16_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_213_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09329_ _18548_/Q _18547_/Q _18546_/Q vssd1 vssd1 vccd1 vccd1 _09332_/B sky130_fd_sc_hd__or3_2
XFILLER_51_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12340_ _12340_/A _12340_/B _12340_/C vssd1 vssd1 vccd1 vccd1 _12340_/X sky130_fd_sc_hd__and3_1
XFILLER_166_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_216_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12271_ _12289_/A vssd1 vssd1 vccd1 vccd1 _12304_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_119_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14010_ _11957_/B _13875_/X _13924_/X _14009_/X vssd1 vssd1 vccd1 vccd1 _14010_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_153_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11222_ _11224_/A _11224_/C _11221_/X vssd1 vssd1 vccd1 vccd1 _11222_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_4_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19103__74 vssd1 vssd1 vccd1 vccd1 _19103__74/HI _19211_/A sky130_fd_sc_hd__conb_1
XFILLER_218_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11153_ _11584_/B vssd1 vssd1 vccd1 vccd1 _11770_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_122_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10104_ _09260_/B _10060_/X _10103_/X _09987_/A vssd1 vssd1 vccd1 vccd1 _10104_/X
+ sky130_fd_sc_hd__o211a_1
X_15961_ _15960_/B _15956_/X _15960_/Y _15948_/X vssd1 vssd1 vccd1 vccd1 _18566_/D
+ sky130_fd_sc_hd__o211a_1
X_11084_ _17791_/Q vssd1 vssd1 vccd1 vccd1 _11951_/A sky130_fd_sc_hd__buf_2
XFILLER_62_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14912_ _18353_/Q _18317_/Q _14934_/S vssd1 vssd1 vccd1 vccd1 _14912_/X sky130_fd_sc_hd__mux2_1
X_10035_ _09198_/A _09193_/A _09203_/B _10293_/A _10025_/A _09986_/A vssd1 vssd1 vccd1
+ vccd1 _10035_/X sky130_fd_sc_hd__mux4_1
X_17700_ _17700_/A vssd1 vssd1 vccd1 vccd1 _18987_/D sky130_fd_sc_hd__clkbuf_1
XTAP_5464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18680_ _18682_/CLK _18680_/D vssd1 vssd1 vccd1 vccd1 _18680_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_209_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15892_ _16041_/A _15892_/B vssd1 vssd1 vccd1 vccd1 _15900_/B sky130_fd_sc_hd__nor2_2
XTAP_4730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14843_ _14856_/A _15279_/B _14843_/C vssd1 vssd1 vccd1 vccd1 _14843_/X sky130_fd_sc_hd__or3_1
X_17631_ _17631_/A vssd1 vssd1 vccd1 vccd1 _17631_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_84_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17562_ _17560_/Y _17552_/A _14414_/A vssd1 vssd1 vccd1 vccd1 _17562_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_84_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14774_ _18282_/Q _14777_/B _14773_/X _14758_/X vssd1 vssd1 vccd1 vccd1 _18282_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_95_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11986_ _11963_/A _11944_/A _11976_/A _11932_/A vssd1 vssd1 vccd1 vccd1 _11988_/C
+ sky130_fd_sc_hd__a22o_1
X_16513_ _17120_/A _16976_/B vssd1 vssd1 vccd1 vccd1 _16578_/A sky130_fd_sc_hd__or2_2
XFILLER_186_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13725_ _13743_/A vssd1 vssd1 vccd1 vccd1 _13725_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_16_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_186_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17493_ _17493_/A _17493_/B _17516_/C vssd1 vssd1 vccd1 vccd1 _17493_/X sky130_fd_sc_hd__or3_1
X_10937_ _10547_/B _10930_/X _10936_/X _10512_/B vssd1 vssd1 vccd1 vccd1 _10937_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_205_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_204_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_220_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16444_ _16491_/A _16736_/B _16481_/C vssd1 vssd1 vccd1 vccd1 _16444_/X sky130_fd_sc_hd__or3_1
XFILLER_143_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19232_ _19232_/A _08937_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[32] sky130_fd_sc_hd__ebufn_8
XFILLER_31_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13656_ _18963_/Q _13654_/X _13592_/A _18978_/Q _13655_/X vssd1 vssd1 vccd1 vccd1
+ _13656_/X sky130_fd_sc_hd__a221o_1
XFILLER_108_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10868_ _14247_/A _10865_/X _10867_/X _10843_/X vssd1 vssd1 vccd1 vccd1 _10868_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_176_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_176_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19163_ _19163_/A _09026_/Y vssd1 vssd1 vccd1 vccd1 io_out[1] sky130_fd_sc_hd__ebufn_8
XFILLER_220_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12607_ _12607_/A vssd1 vssd1 vccd1 vccd1 _12618_/A sky130_fd_sc_hd__inv_2
X_16375_ _16780_/A vssd1 vssd1 vccd1 vccd1 _16456_/A sky130_fd_sc_hd__clkbuf_2
XPHY_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13587_ _13857_/A vssd1 vssd1 vccd1 vccd1 _13588_/A sky130_fd_sc_hd__buf_6
XFILLER_129_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_185_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10799_ _09165_/A _09160_/C _09170_/D _10308_/A _10770_/A _10781_/S vssd1 vssd1 vccd1
+ vccd1 _10799_/X sky130_fd_sc_hd__mux4_1
XFILLER_9_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18114_ _18114_/CLK _18114_/D vssd1 vssd1 vccd1 vccd1 _18114_/Q sky130_fd_sc_hd__dfxtp_1
X_15326_ _15325_/B _15322_/X _15325_/Y _15315_/X vssd1 vssd1 vccd1 vccd1 _18416_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_184_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12538_ _14185_/A _12538_/B vssd1 vssd1 vccd1 vccd1 _17917_/D sky130_fd_sc_hd__nand2_1
XFILLER_145_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18045_ _18052_/CLK _18045_/D vssd1 vssd1 vccd1 vccd1 _18045_/Q sky130_fd_sc_hd__dfxtp_1
X_15257_ _15279_/A _15257_/B _15257_/C vssd1 vssd1 vccd1 vccd1 _15257_/X sky130_fd_sc_hd__or3_1
XFILLER_172_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_126_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12469_ _17905_/Q _12487_/B _12465_/Y vssd1 vssd1 vccd1 vccd1 _12471_/A sky130_fd_sc_hd__a21o_1
X_14208_ _14207_/X _09935_/X _14267_/A vssd1 vssd1 vccd1 vccd1 _14208_/X sky130_fd_sc_hd__mux2_1
X_15188_ _15195_/B _15185_/X _15186_/X _15187_/X vssd1 vssd1 vccd1 vccd1 _18384_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_158_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14139_ _18365_/Q _13697_/A _13537_/A _18341_/Q vssd1 vssd1 vccd1 vccd1 _14139_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_67_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18947_ _18953_/CLK _18947_/D vssd1 vssd1 vccd1 vccd1 _18947_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_101_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_1344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_228_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09680_ _12078_/A _09699_/B vssd1 vssd1 vccd1 vccd1 _10046_/A sky130_fd_sc_hd__xor2_4
XFILLER_66_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18878_ _18914_/CLK _18878_/D vssd1 vssd1 vccd1 vccd1 _18878_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_95_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_143_wb_clk_i clkbuf_5_26_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18290_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_17829_ _18209_/CLK _17829_/D vssd1 vssd1 vccd1 vccd1 _17829_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_81_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_222_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_206_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09114_ _09114_/A _09114_/B _09114_/C _10728_/A vssd1 vssd1 vccd1 vccd1 _09120_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_182_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09045_ _09046_/A vssd1 vssd1 vccd1 vccd1 _09045_/Y sky130_fd_sc_hd__inv_2
XFILLER_190_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_163_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_164_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_1282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_5_14_0_wb_clk_i clkbuf_4_7_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18114_/CLK
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_104_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09947_ _09947_/A vssd1 vssd1 vccd1 vccd1 _09948_/A sky130_fd_sc_hd__buf_2
XFILLER_104_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_213_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_10 _09148_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_21 _09214_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09878_ _09901_/A _09907_/A vssd1 vssd1 vccd1 vccd1 _09902_/A sky130_fd_sc_hd__nor2_4
XTAP_4037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_32 _09688_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_43 _10068_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_54 _15840_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_65 _13763_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_76 _13538_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_87 _13625_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_98 _13781_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11840_ _11526_/B _11528_/X _11848_/A vssd1 vssd1 vccd1 vccd1 _11840_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_2_1344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11771_ _11770_/A _11770_/C _11770_/B vssd1 vssd1 vccd1 vccd1 _11772_/B sky130_fd_sc_hd__a21oi_1
XTAP_1934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13510_ _13563_/A _13557_/B vssd1 vssd1 vccd1 vccd1 _13667_/A sky130_fd_sc_hd__nor2_2
XFILLER_14_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10722_ _10722_/A _10763_/S vssd1 vssd1 vccd1 vccd1 _10722_/X sky130_fd_sc_hd__or2_1
XTAP_1967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14490_ _14490_/A vssd1 vssd1 vccd1 vccd1 _18219_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13441_ _11070_/X _13422_/Y _13426_/Y vssd1 vssd1 vccd1 vccd1 _13441_/X sky130_fd_sc_hd__a21o_1
XFILLER_201_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10653_ _10689_/A vssd1 vssd1 vccd1 vccd1 _10867_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_201_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16160_ _16202_/A _16160_/B vssd1 vssd1 vccd1 vccd1 _16160_/Y sky130_fd_sc_hd__nand2_1
XFILLER_10_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13372_ _13372_/A _13389_/B vssd1 vssd1 vccd1 vccd1 _13372_/Y sky130_fd_sc_hd__nand2_1
X_10584_ _10582_/S _10583_/X _10029_/S vssd1 vssd1 vccd1 vccd1 _10584_/X sky130_fd_sc_hd__a21o_1
XFILLER_220_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15111_ _15232_/A vssd1 vssd1 vccd1 vccd1 _15162_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_127_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12323_ _12323_/A _12323_/B _12323_/C vssd1 vssd1 vccd1 vccd1 _12323_/X sky130_fd_sc_hd__and3_1
X_16091_ _18634_/Q _18598_/Q _16091_/S vssd1 vssd1 vccd1 vccd1 _16091_/X sky130_fd_sc_hd__mux2_1
XFILLER_181_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15042_ _15042_/A _15186_/B _15054_/C vssd1 vssd1 vccd1 vccd1 _15042_/X sky130_fd_sc_hd__or3_1
XFILLER_119_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12254_ _12269_/B _12269_/C vssd1 vssd1 vccd1 vccd1 _12270_/A sky130_fd_sc_hd__nand2_1
XFILLER_123_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11205_ _17813_/Q _17812_/Q _11205_/C vssd1 vssd1 vccd1 vccd1 _11209_/B sky130_fd_sc_hd__nand3_1
XFILLER_64_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12185_ _12180_/Y _12183_/X _12184_/X vssd1 vssd1 vccd1 vccd1 _17849_/D sky130_fd_sc_hd__o21a_1
X_18801_ _18806_/CLK _18801_/D vssd1 vssd1 vccd1 vccd1 _18801_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_96_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11136_ _11661_/A vssd1 vssd1 vccd1 vccd1 _11253_/A sky130_fd_sc_hd__buf_2
XFILLER_190_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16993_ _16998_/B _16991_/X _16992_/X _16964_/X vssd1 vssd1 vccd1 vccd1 _18810_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_27_1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18732_ _18732_/CLK _18732_/D vssd1 vssd1 vccd1 vccd1 _18732_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_62_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15944_ _15944_/A _15993_/B vssd1 vssd1 vccd1 vccd1 _15960_/B sky130_fd_sc_hd__nor2_2
XTAP_5250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11067_ _11970_/C vssd1 vssd1 vccd1 vccd1 _11334_/B sky130_fd_sc_hd__clkbuf_2
XTAP_5261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10018_ _09119_/C _09109_/C _10019_/S vssd1 vssd1 vccd1 vccd1 _10018_/X sky130_fd_sc_hd__mux2_1
XTAP_5294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18663_ _18663_/CLK _18663_/D vssd1 vssd1 vccd1 vccd1 _18663_/Q sky130_fd_sc_hd__dfxtp_1
X_15875_ _18584_/Q _18548_/Q _15879_/S vssd1 vssd1 vccd1 vccd1 _15875_/X sky130_fd_sc_hd__mux2_1
XFILLER_37_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_221_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14826_ _14948_/A vssd1 vssd1 vccd1 vccd1 _14875_/A sky130_fd_sc_hd__clkbuf_2
X_17614_ _17638_/A _17614_/B vssd1 vssd1 vccd1 vccd1 _17615_/A sky130_fd_sc_hd__and2_1
XFILLER_92_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18594_ _18633_/CLK _18594_/D vssd1 vssd1 vccd1 vccd1 _18594_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_3870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14757_ _14793_/A _15199_/B _14757_/C vssd1 vssd1 vccd1 vccd1 _14757_/X sky130_fd_sc_hd__or3_1
X_17545_ _17544_/B _17543_/X _17544_/Y _11816_/X vssd1 vssd1 vccd1 vccd1 _18950_/D
+ sky130_fd_sc_hd__o211a_1
X_11969_ _11948_/X _11946_/X _11968_/X _11973_/A vssd1 vssd1 vccd1 vccd1 _12022_/A
+ sky130_fd_sc_hd__a211oi_1
X_13708_ _18750_/Q _13834_/A _13704_/X _13707_/X vssd1 vssd1 vccd1 vccd1 _13708_/X
+ sky130_fd_sc_hd__a211o_1
X_17476_ _18931_/Q _17477_/B _17475_/Y _17461_/X vssd1 vssd1 vccd1 vccd1 _18931_/D
+ sky130_fd_sc_hd__o211a_1
X_14688_ _16959_/A vssd1 vssd1 vccd1 vccd1 _16962_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_32_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19215_ _19215_/A _08968_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[15] sky130_fd_sc_hd__ebufn_8
X_16427_ _16429_/B _16425_/X _16426_/Y _16418_/X vssd1 vssd1 vccd1 vccd1 _18676_/D
+ sky130_fd_sc_hd__o211a_1
X_13639_ _18894_/Q _13702_/A _13625_/X _18888_/Q _13638_/X vssd1 vssd1 vccd1 vccd1
+ _13639_/X sky130_fd_sc_hd__a221o_1
XFILLER_220_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16358_ _16371_/A _16796_/B _16358_/C vssd1 vssd1 vccd1 vccd1 _16358_/X sky130_fd_sc_hd__or3_1
X_19146_ _19146_/A _09045_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[16] sky130_fd_sc_hd__ebufn_8
XFILLER_185_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_1176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15309_ _15415_/A vssd1 vssd1 vccd1 vccd1 _15334_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_69_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_157_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16289_ _16289_/A vssd1 vssd1 vccd1 vccd1 _16333_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_195_1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18028_ _18087_/CLK _18028_/D vssd1 vssd1 vccd1 vccd1 _18028_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_133_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09801_ _09752_/A _09746_/B _09800_/X vssd1 vssd1 vccd1 vccd1 _09807_/A sky130_fd_sc_hd__a21o_1
XFILLER_113_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19094__65 vssd1 vssd1 vccd1 vccd1 _19094__65/HI _19202_/A sky130_fd_sc_hd__conb_1
XFILLER_45_1272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09732_ _09742_/A _09732_/B vssd1 vssd1 vccd1 vccd1 _09739_/B sky130_fd_sc_hd__xnor2_1
XFILLER_86_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_228_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_189_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_189_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19129__100 vssd1 vssd1 vccd1 vccd1 _19129__100/HI _19237_/A sky130_fd_sc_hd__conb_1
X_09663_ _12079_/A _12080_/S vssd1 vssd1 vccd1 vccd1 _09664_/B sky130_fd_sc_hd__xnor2_1
XFILLER_54_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_215_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_1316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09594_ _09593_/A _09593_/B _09593_/C vssd1 vssd1 vccd1 vccd1 _09594_/X sky130_fd_sc_hd__o21a_1
XFILLER_215_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_231_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINSDIODE2_180 _08954_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_210_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_191 _09119_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_210_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_40_wb_clk_i _18759_/CLK vssd1 vssd1 vccd1 vccd1 _18765_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_149_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09028_ _09028_/A vssd1 vssd1 vccd1 vccd1 _09028_/Y sky130_fd_sc_hd__inv_2
XFILLER_191_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_105_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13990_ _18409_/Q _13758_/A _13841_/A _18385_/Q _13989_/X vssd1 vssd1 vccd1 vccd1
+ _13990_/X sky130_fd_sc_hd__a221o_1
XFILLER_77_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_218_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_213_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12941_ _11036_/B _12951_/A _12930_/A vssd1 vssd1 vccd1 vccd1 _12941_/Y sky130_fd_sc_hd__o21ai_1
XTAP_3100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_218_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15660_ _18530_/Q _18494_/Q _15665_/S vssd1 vssd1 vccd1 vccd1 _15660_/X sky130_fd_sc_hd__mux2_1
XTAP_3144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12872_ _17954_/Q _12869_/A _12862_/X vssd1 vssd1 vccd1 vccd1 _12873_/B sky130_fd_sc_hd__o21ai_1
XTAP_2410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14611_ _17471_/A vssd1 vssd1 vccd1 vccd1 _14612_/A sky130_fd_sc_hd__buf_2
XFILLER_27_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11823_ _18155_/Q _11813_/Y _11820_/X _11717_/Y _11822_/X vssd1 vssd1 vccd1 vccd1
+ _17826_/D sky130_fd_sc_hd__o221a_1
XFILLER_61_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15591_ _15630_/A _15594_/B vssd1 vssd1 vccd1 vccd1 _15591_/Y sky130_fd_sc_hd__nand2_1
XTAP_1720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17330_ _17448_/A vssd1 vssd1 vccd1 vccd1 _17376_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_199_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14542_ _15957_/A vssd1 vssd1 vccd1 vccd1 _15649_/A sky130_fd_sc_hd__buf_12
XFILLER_121_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11754_ _17915_/Q vssd1 vssd1 vccd1 vccd1 _11767_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_109_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10705_ _10705_/A vssd1 vssd1 vccd1 vccd1 _13000_/A sky130_fd_sc_hd__clkbuf_4
X_17261_ _17263_/B _17258_/X _17259_/Y _17260_/X vssd1 vssd1 vccd1 vccd1 _18877_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_187_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14473_ _14214_/Y _14471_/C _17766_/A vssd1 vssd1 vccd1 vccd1 _18211_/D sky130_fd_sc_hd__a21oi_1
X_11685_ _17853_/Q vssd1 vssd1 vccd1 vccd1 _11685_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_16212_ _16212_/A vssd1 vssd1 vccd1 vccd1 _16265_/A sky130_fd_sc_hd__buf_2
X_19000_ _19000_/CLK _19000_/D vssd1 vssd1 vccd1 vccd1 _19000_/Q sky130_fd_sc_hd__dfxtp_1
X_13424_ _13648_/A _13649_/B vssd1 vssd1 vccd1 vccd1 _13435_/B sky130_fd_sc_hd__nand2_1
XFILLER_14_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10636_ _12074_/A _12966_/A _10650_/B vssd1 vssd1 vccd1 vccd1 _12096_/B sky130_fd_sc_hd__and3_2
X_17192_ _18897_/Q _18861_/Q _17199_/S vssd1 vssd1 vccd1 vccd1 _17192_/X sky130_fd_sc_hd__mux2_1
X_16143_ _16199_/A _16147_/B vssd1 vssd1 vccd1 vccd1 _16143_/Y sky130_fd_sc_hd__nand2_1
X_13355_ _17779_/Q _17780_/Q vssd1 vssd1 vccd1 vccd1 _13356_/B sky130_fd_sc_hd__or2_1
XFILLER_182_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10567_ _09294_/A _09304_/B _10575_/B vssd1 vssd1 vccd1 vccd1 _10567_/X sky130_fd_sc_hd__mux2_1
XFILLER_155_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_154_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12306_ _12327_/A _12327_/B vssd1 vssd1 vccd1 vccd1 _12329_/C sky130_fd_sc_hd__and2_1
X_16074_ _16139_/A vssd1 vssd1 vccd1 vccd1 _16074_/X sky130_fd_sc_hd__clkbuf_2
X_13286_ _13286_/A _13286_/B _13286_/C _13286_/D vssd1 vssd1 vccd1 vccd1 _13292_/C
+ sky130_fd_sc_hd__or4_1
XFILLER_154_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10498_ _10498_/A _10497_/X vssd1 vssd1 vccd1 vccd1 _10498_/X sky130_fd_sc_hd__or2b_2
XFILLER_143_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_170_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15025_ _15061_/A _15025_/B vssd1 vssd1 vccd1 vccd1 _15025_/Y sky130_fd_sc_hd__nand2_1
XFILLER_68_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_216_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12237_ _12246_/A vssd1 vssd1 vccd1 vccd1 _12258_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_190_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12168_ _12169_/A _12169_/B vssd1 vssd1 vccd1 vccd1 _12168_/X sky130_fd_sc_hd__and2_1
XFILLER_2_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11119_ _11735_/A vssd1 vssd1 vccd1 vccd1 _11748_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_96_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16976_ _17549_/A _16976_/B vssd1 vssd1 vccd1 vccd1 _17012_/A sky130_fd_sc_hd__or2_1
X_12099_ _12099_/A _12099_/B vssd1 vssd1 vccd1 vccd1 _12103_/A sky130_fd_sc_hd__xnor2_1
XFILLER_7_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18715_ _18719_/CLK _18715_/D vssd1 vssd1 vccd1 vccd1 _18715_/Q sky130_fd_sc_hd__dfxtp_2
X_15927_ _18596_/Q _18560_/Q _15937_/S vssd1 vssd1 vccd1 vccd1 _15927_/X sky130_fd_sc_hd__mux2_1
XTAP_5080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput6 io_in[28] vssd1 vssd1 vccd1 vccd1 input6/X sky130_fd_sc_hd__clkbuf_1
XTAP_5091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18646_ _18682_/CLK _18646_/D vssd1 vssd1 vccd1 vccd1 _18646_/Q sky130_fd_sc_hd__dfxtp_2
X_15858_ _15865_/B _15856_/X _15857_/X _15842_/X vssd1 vssd1 vccd1 vccd1 _18543_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_4390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14809_ _18328_/Q _18292_/Q _14809_/S vssd1 vssd1 vccd1 vccd1 _14809_/X sky130_fd_sc_hd__mux2_1
XFILLER_91_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_206_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18577_ _18577_/CLK _18577_/D vssd1 vssd1 vccd1 vccd1 _18577_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_18_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15789_ _15795_/B _15787_/X _15788_/X _15783_/X vssd1 vssd1 vccd1 vccd1 _18525_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_33_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17528_ _17538_/A _17528_/B _17538_/C vssd1 vssd1 vccd1 vccd1 _17528_/X sky130_fd_sc_hd__or3_1
XFILLER_189_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_1208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17459_ _18963_/Q _18927_/Q _17467_/S vssd1 vssd1 vccd1 vccd1 _17459_/X sky130_fd_sc_hd__mux2_1
XFILLER_193_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_221_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_192_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_214_1350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09715_ _18260_/Q _18259_/Q _18258_/Q vssd1 vssd1 vccd1 vccd1 _09715_/X sky130_fd_sc_hd__or3_4
XFILLER_19_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09646_ _09647_/A _09647_/B vssd1 vssd1 vccd1 vccd1 _09649_/B sky130_fd_sc_hd__nor2_1
XFILLER_16_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_222_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_204_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09577_ _18108_/Q _17981_/Q vssd1 vssd1 vccd1 vccd1 _09578_/B sky130_fd_sc_hd__xnor2_1
XTAP_1027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_208_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_212_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11470_ _11482_/A _11482_/B _11483_/B vssd1 vssd1 vccd1 vccd1 _11470_/Y sky130_fd_sc_hd__nor3b_1
XFILLER_11_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_221_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_183_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10421_ _10419_/A _10420_/X _10918_/S vssd1 vssd1 vccd1 vccd1 _10421_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_104_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13140_ _13140_/A _18030_/Q vssd1 vssd1 vccd1 vccd1 _13141_/A sky130_fd_sc_hd__and2_1
X_10352_ _14240_/B _10349_/X _10351_/X _10388_/A vssd1 vssd1 vccd1 vccd1 _10352_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_192_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_100_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_174_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13071_ _13071_/A vssd1 vssd1 vccd1 vccd1 _18000_/D sky130_fd_sc_hd__clkbuf_1
X_10283_ _09176_/A _09186_/D _12123_/A vssd1 vssd1 vccd1 vccd1 _10283_/X sky130_fd_sc_hd__mux2_1
XFILLER_183_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12022_ _12022_/A _12022_/B _12022_/C _12042_/A vssd1 vssd1 vccd1 vccd1 _12028_/B
+ sky130_fd_sc_hd__or4_1
XFILLER_105_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_215_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16830_ _16833_/B _16827_/X _16829_/Y _16825_/X vssd1 vssd1 vccd1 vccd1 _18775_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_78_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16761_ _16769_/B _16758_/X _16759_/X _16760_/X vssd1 vssd1 vccd1 vccd1 _18759_/D
+ sky130_fd_sc_hd__o211a_1
X_13973_ _18271_/Q _13735_/X _13764_/X _18295_/Q vssd1 vssd1 vccd1 vccd1 _13973_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_24_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18500_ _18504_/CLK _18500_/D vssd1 vssd1 vccd1 vccd1 _18500_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_4_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15712_ _15734_/A _16007_/B _15724_/C vssd1 vssd1 vccd1 vccd1 _15712_/X sky130_fd_sc_hd__or3_1
XFILLER_185_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12924_ _13318_/A _12924_/B vssd1 vssd1 vccd1 vccd1 _12924_/Y sky130_fd_sc_hd__nor2_1
X_16692_ _16736_/A _16692_/B _16716_/C vssd1 vssd1 vccd1 vccd1 _16692_/X sky130_fd_sc_hd__or3_1
XFILLER_19_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_1216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_5_7_0_wb_clk_i clkbuf_5_7_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_5_7_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_185_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18431_ _18432_/CLK _18431_/D vssd1 vssd1 vccd1 vccd1 _18431_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_59_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_1298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15643_ _15643_/A vssd1 vssd1 vccd1 vccd1 _15885_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_185_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12855_ _12816_/X _12857_/C _12854_/X vssd1 vssd1 vccd1 vccd1 _12855_/Y sky130_fd_sc_hd__o21ai_1
XTAP_2240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11806_ _11970_/C _11806_/B vssd1 vssd1 vccd1 vccd1 _11937_/C sky130_fd_sc_hd__or2_2
X_15574_ _15613_/A _16021_/B _15574_/C vssd1 vssd1 vccd1 vccd1 _15574_/X sky130_fd_sc_hd__or3_1
X_18362_ _18393_/CLK _18362_/D vssd1 vssd1 vccd1 vccd1 _18362_/Q sky130_fd_sc_hd__dfxtp_4
XTAP_2284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12786_ _17943_/Q _12786_/B vssd1 vssd1 vccd1 vccd1 _12786_/X sky130_fd_sc_hd__or2_1
XTAP_2295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14525_ _16512_/C _15463_/B _15607_/B _15903_/C vssd1 vssd1 vccd1 vccd1 _14526_/B
+ sky130_fd_sc_hd__or4b_1
X_17313_ _18926_/Q _18890_/Q _17317_/S vssd1 vssd1 vccd1 vccd1 _17313_/X sky130_fd_sc_hd__mux2_1
XFILLER_159_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11737_ _17914_/Q _11737_/B vssd1 vssd1 vccd1 vccd1 _11760_/B sky130_fd_sc_hd__and2_1
XFILLER_109_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18293_ _18312_/CLK _18293_/D vssd1 vssd1 vccd1 vccd1 _18293_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_187_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17244_ _18909_/Q _18873_/Q _17244_/S vssd1 vssd1 vccd1 vccd1 _17244_/X sky130_fd_sc_hd__mux2_1
XFILLER_30_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14456_ _14404_/X _09506_/B _14405_/X vssd1 vssd1 vccd1 vccd1 _14457_/C sky130_fd_sc_hd__a21o_1
XFILLER_70_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11668_ _11668_/A _11668_/B vssd1 vssd1 vccd1 vccd1 _11669_/C sky130_fd_sc_hd__nor2_1
XFILLER_186_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13407_ _18129_/Q _11040_/X _11035_/B _13381_/X _13395_/X vssd1 vssd1 vccd1 vccd1
+ _18129_/D sky130_fd_sc_hd__o2111a_1
X_10619_ _10619_/A _10619_/B vssd1 vssd1 vccd1 vccd1 _10619_/Y sky130_fd_sc_hd__nor2_1
X_17175_ _17226_/A vssd1 vssd1 vccd1 vccd1 _17199_/S sky130_fd_sc_hd__clkbuf_2
X_14387_ _18189_/Q _14384_/A _14384_/B _12972_/A vssd1 vssd1 vccd1 vccd1 _14387_/X
+ sky130_fd_sc_hd__a31o_1
X_11599_ _17858_/Q vssd1 vssd1 vccd1 vccd1 _11603_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_116_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16126_ _16193_/A vssd1 vssd1 vccd1 vccd1 _16181_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_196_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13338_ _13375_/A _13394_/D _13375_/B _13375_/C vssd1 vssd1 vccd1 vccd1 _17768_/B
+ sky130_fd_sc_hd__nor4_4
XFILLER_192_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16057_ _16219_/A vssd1 vssd1 vccd1 vccd1 _16666_/B sky130_fd_sc_hd__buf_4
X_13269_ _18153_/Q _13269_/B vssd1 vssd1 vccd1 vccd1 _13269_/X sky130_fd_sc_hd__or2_1
XFILLER_44_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15008_ _15058_/A _15012_/B vssd1 vssd1 vccd1 vccd1 _15008_/Y sky130_fd_sc_hd__nand2_1
XFILLER_102_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_97_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19064__35 vssd1 vssd1 vccd1 vccd1 _19064__35/HI _19158_/A sky130_fd_sc_hd__conb_1
XFILLER_96_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16959_ _16959_/A vssd1 vssd1 vccd1 vccd1 _17536_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_2_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09500_ _18198_/Q _09500_/B vssd1 vssd1 vccd1 vccd1 _09501_/B sky130_fd_sc_hd__or2_1
XFILLER_110_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09431_ _09431_/A vssd1 vssd1 vccd1 vccd1 _09432_/B sky130_fd_sc_hd__inv_2
XFILLER_65_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_227_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18629_ _18650_/CLK _18629_/D vssd1 vssd1 vccd1 vccd1 _18629_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_80_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09362_ _18293_/Q _18292_/Q _18291_/Q vssd1 vssd1 vccd1 vccd1 _09365_/B sky130_fd_sc_hd__or3_4
XFILLER_40_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_221_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09293_ _18494_/Q _18493_/Q _18492_/Q vssd1 vssd1 vccd1 vccd1 _09294_/D sky130_fd_sc_hd__or3_4
XFILLER_20_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_178_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_217_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_142_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_210_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10970_ _18228_/Q vssd1 vssd1 vccd1 vccd1 _14515_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_216_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_210_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09629_ _09665_/A _09665_/B vssd1 vssd1 vccd1 vccd1 _09630_/B sky130_fd_sc_hd__xnor2_4
XFILLER_16_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12640_ _12640_/A _12640_/B vssd1 vssd1 vccd1 vccd1 _12640_/Y sky130_fd_sc_hd__nand2_1
XFILLER_31_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_203_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12571_ _12556_/A _12564_/X _12556_/B _12570_/Y _12554_/B vssd1 vssd1 vccd1 vccd1
+ _12571_/X sky130_fd_sc_hd__a311o_2
XFILLER_169_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_1274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14310_ _14311_/A _14311_/B vssd1 vssd1 vccd1 vccd1 _14310_/Y sky130_fd_sc_hd__nor2_1
X_11522_ _11522_/A _12285_/B _12285_/C vssd1 vssd1 vccd1 vccd1 _11522_/X sky130_fd_sc_hd__and3_1
X_15290_ _17120_/A _15757_/A vssd1 vssd1 vccd1 vccd1 _15370_/A sky130_fd_sc_hd__or2_2
XFILLER_178_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_211_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_184_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14241_ _14260_/A _14239_/Y _14240_/Y _14272_/A vssd1 vssd1 vccd1 vccd1 _14241_/X
+ sky130_fd_sc_hd__o211a_1
X_11453_ _11453_/A _11453_/B vssd1 vssd1 vccd1 vccd1 _11482_/A sky130_fd_sc_hd__xor2_1
X_10404_ _10399_/X _10403_/X _09889_/X vssd1 vssd1 vccd1 vccd1 _10404_/Y sky130_fd_sc_hd__a21boi_1
XFILLER_109_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14172_ _18623_/Q _13838_/A _14170_/X _14171_/X vssd1 vssd1 vccd1 vccd1 _14172_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_165_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_137_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11384_ _11384_/A vssd1 vssd1 vccd1 vccd1 _11384_/Y sky130_fd_sc_hd__inv_2
XFILLER_152_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_109_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_194_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13123_ _13129_/A _18022_/Q vssd1 vssd1 vccd1 vccd1 _13124_/A sky130_fd_sc_hd__and2_1
XFILLER_98_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10335_ _10338_/A _09889_/X _10329_/X _10334_/X _09930_/X vssd1 vssd1 vccd1 vccd1
+ _10335_/X sky130_fd_sc_hd__a32o_1
XFILLER_11_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18980_ _18980_/CLK _18980_/D vssd1 vssd1 vccd1 vccd1 _18980_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_180_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13054_ _13052_/X _13055_/B _18002_/Q vssd1 vssd1 vccd1 vccd1 _13054_/Y sky130_fd_sc_hd__o21ai_1
X_17931_ _17931_/CLK _17931_/D vssd1 vssd1 vccd1 vccd1 _17931_/Q sky130_fd_sc_hd__dfxtp_1
X_10266_ _11924_/A _10237_/X _10265_/X vssd1 vssd1 vccd1 vccd1 _10270_/B sky130_fd_sc_hd__a21o_1
XFILLER_105_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12005_ _12025_/B _11946_/X _12004_/Y _11948_/X vssd1 vssd1 vccd1 vccd1 _12018_/A
+ sky130_fd_sc_hd__a31o_2
XFILLER_6_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17862_ _19035_/CLK _17862_/D vssd1 vssd1 vccd1 vccd1 _17862_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_65_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10197_ _10197_/A _10197_/B vssd1 vssd1 vccd1 vccd1 _10201_/B sky130_fd_sc_hd__xnor2_1
XFILLER_121_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16813_ _16813_/A _16815_/B vssd1 vssd1 vccd1 vccd1 _16813_/Y sky130_fd_sc_hd__nand2_1
XFILLER_93_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17793_ _17793_/CLK _17793_/D vssd1 vssd1 vccd1 vccd1 _17793_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_94_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16744_ _16743_/B _16742_/X _16743_/Y _16740_/X vssd1 vssd1 vccd1 vccd1 _18755_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_81_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13956_ _18643_/Q _13772_/X _13752_/X _18637_/Q vssd1 vssd1 vccd1 vccd1 _13956_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_4_1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12907_ _12907_/A vssd1 vssd1 vccd1 vccd1 _17965_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_207_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16675_ _16787_/A vssd1 vssd1 vccd1 vccd1 _16766_/A sky130_fd_sc_hd__buf_2
X_13887_ _18970_/Q _13705_/A _13706_/A _18952_/Q vssd1 vssd1 vccd1 vccd1 _13887_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_228_1338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_222_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_185_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18414_ _18416_/CLK _18414_/D vssd1 vssd1 vccd1 vccd1 _18414_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_146_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15626_ _15869_/A vssd1 vssd1 vccd1 vccd1 _15678_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_34_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12838_ _12874_/A vssd1 vssd1 vccd1 vccd1 _12888_/B sky130_fd_sc_hd__clkbuf_2
XTAP_2070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_210_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18345_ _18346_/CLK _18345_/D vssd1 vssd1 vccd1 vccd1 _18345_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_124_1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15557_ _18506_/Q _18470_/Q _15565_/S vssd1 vssd1 vccd1 vccd1 _15557_/X sky130_fd_sc_hd__mux2_1
X_12769_ _13318_/B _13318_/C vssd1 vssd1 vccd1 vccd1 _12769_/Y sky130_fd_sc_hd__nor2_1
XTAP_1380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_159_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_1208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_147_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_168_wb_clk_i clkbuf_5_10_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18030_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_14508_ _14508_/A _14513_/B vssd1 vssd1 vccd1 vccd1 _14515_/C sky130_fd_sc_hd__or2_1
X_15488_ _15487_/B _15486_/X _15487_/Y _15474_/X vssd1 vssd1 vccd1 vccd1 _18452_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_187_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18276_ _18278_/CLK _18276_/D vssd1 vssd1 vccd1 vccd1 _18276_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_124_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19109__80 vssd1 vssd1 vccd1 vccd1 _19109__80/HI _19217_/A sky130_fd_sc_hd__conb_1
X_17227_ _18905_/Q _18869_/Q _17244_/S vssd1 vssd1 vccd1 vccd1 _17227_/X sky130_fd_sc_hd__mux2_1
X_14439_ _09503_/B _14428_/A _14434_/Y _14438_/Y vssd1 vssd1 vccd1 vccd1 _14440_/B
+ sky130_fd_sc_hd__o22ai_1
XFILLER_190_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17158_ _17446_/A _17202_/B vssd1 vssd1 vccd1 vccd1 _17169_/B sky130_fd_sc_hd__nor2_2
XFILLER_171_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16109_ _16132_/A _16109_/B vssd1 vssd1 vccd1 vccd1 _16109_/Y sky130_fd_sc_hd__nand2_1
XFILLER_196_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17089_ _17091_/B _17087_/X _17088_/Y _17076_/X vssd1 vssd1 vccd1 vccd1 _18835_/D
+ sky130_fd_sc_hd__o211a_1
X_09980_ _12126_/A vssd1 vssd1 vccd1 vccd1 _09981_/A sky130_fd_sc_hd__buf_2
XFILLER_131_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_1331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08931_ _08935_/A vssd1 vssd1 vccd1 vccd1 _08931_/Y sky130_fd_sc_hd__inv_2
XFILLER_157_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_229_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_229_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_1307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_226_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_226_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_225_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09414_ _18314_/Q _18313_/Q _18312_/Q vssd1 vssd1 vccd1 vccd1 _09418_/A sky130_fd_sc_hd__or3_1
XFILLER_13_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09345_ _18440_/Q _18439_/Q _18438_/Q vssd1 vssd1 vccd1 vccd1 _09349_/A sky130_fd_sc_hd__or3_4
XFILLER_205_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_178_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09276_ _18878_/Q _18877_/Q _18876_/Q vssd1 vssd1 vccd1 vccd1 _09277_/D sky130_fd_sc_hd__or3_2
XFILLER_138_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_161_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10120_ _10120_/A _10120_/B _10120_/C vssd1 vssd1 vccd1 vccd1 _10121_/B sky130_fd_sc_hd__and3_1
XFILLER_161_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_216_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10051_ _09203_/A _09198_/C _09193_/D _09203_/D _09682_/A _10019_/S vssd1 vssd1 vccd1
+ vccd1 _10051_/X sky130_fd_sc_hd__mux4_2
XTAP_5624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_216_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13810_ _18381_/Q _13733_/A _13806_/X _13809_/X vssd1 vssd1 vccd1 vccd1 _13810_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_112_1240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14790_ _15229_/A _14790_/B vssd1 vssd1 vccd1 vccd1 _14802_/B sky130_fd_sc_hd__nor2_1
XFILLER_60_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_186_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13741_ _13741_/A vssd1 vssd1 vccd1 vccd1 _13785_/A sky130_fd_sc_hd__buf_4
XFILLER_217_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10953_ _09694_/A _10950_/X _10952_/X _10069_/X vssd1 vssd1 vccd1 vccd1 _10953_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_204_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_217_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_182_1216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_1268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16460_ _16507_/A _16464_/B vssd1 vssd1 vccd1 vccd1 _16460_/Y sky130_fd_sc_hd__nand2_1
X_13672_ _18867_/Q _13670_/X _13766_/A _18843_/Q vssd1 vssd1 vccd1 vccd1 _13672_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_32_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_231_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10884_ _09360_/C _10851_/A _10883_/X _10824_/A vssd1 vssd1 vccd1 vccd1 _10884_/X
+ sky130_fd_sc_hd__o211a_1
XPHY_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15411_ _15417_/B _15408_/X _15410_/X _15404_/X vssd1 vssd1 vccd1 vccd1 _18435_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_188_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12623_ _17927_/Q vssd1 vssd1 vccd1 vccd1 _12627_/B sky130_fd_sc_hd__clkbuf_2
X_16391_ _18704_/Q _18668_/Q _16400_/S vssd1 vssd1 vccd1 vccd1 _16391_/X sky130_fd_sc_hd__mux2_1
XFILLER_31_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_231_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_223_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_145_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15342_ _16853_/A vssd1 vssd1 vccd1 vccd1 _15944_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_212_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_197_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_185_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18130_ _18130_/CLK _18130_/D vssd1 vssd1 vccd1 vccd1 _18130_/Q sky130_fd_sc_hd__dfxtp_2
X_12554_ _12554_/A _12554_/B vssd1 vssd1 vccd1 vccd1 _12557_/A sky130_fd_sc_hd__nor2_1
XFILLER_223_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11505_ _13444_/A _11495_/D _11742_/A _11504_/X vssd1 vssd1 vccd1 vccd1 _11528_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_8_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15273_ _15275_/B _15271_/X _15272_/Y _15264_/X vssd1 vssd1 vccd1 vccd1 _18406_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_32_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18061_ _18061_/CLK _18061_/D vssd1 vssd1 vccd1 vccd1 _18061_/Q sky130_fd_sc_hd__dfxtp_1
X_12485_ _17908_/Q _17907_/Q _12487_/B vssd1 vssd1 vccd1 vccd1 _12485_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_156_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17012_ _17012_/A vssd1 vssd1 vccd1 vccd1 _17070_/B sky130_fd_sc_hd__buf_2
X_14224_ _14279_/A _14305_/A vssd1 vssd1 vccd1 vccd1 _14224_/Y sky130_fd_sc_hd__nand2_1
XFILLER_138_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11436_ _11436_/A vssd1 vssd1 vccd1 vccd1 _11436_/Y sky130_fd_sc_hd__inv_2
XFILLER_32_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14155_ _18755_/Q _14124_/X _13538_/A _18737_/Q vssd1 vssd1 vccd1 vccd1 _14155_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_4_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11367_ _11308_/Y _11577_/B vssd1 vssd1 vccd1 vccd1 _11374_/C sky130_fd_sc_hd__and2b_1
XFILLER_193_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_180_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13106_ _13106_/A vssd1 vssd1 vccd1 vccd1 _18013_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_113_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10318_ _09260_/B _09945_/X _10317_/X _09923_/X vssd1 vssd1 vccd1 vccd1 _10318_/X
+ sky130_fd_sc_hd__o211a_1
X_14086_ _18473_/Q _13532_/A _13539_/A _18449_/Q vssd1 vssd1 vccd1 vccd1 _14086_/X
+ sky130_fd_sc_hd__a22o_1
X_18963_ _18970_/CLK _18963_/D vssd1 vssd1 vccd1 vccd1 _18963_/Q sky130_fd_sc_hd__dfxtp_2
X_11298_ _11297_/B _11297_/C _11313_/B vssd1 vssd1 vccd1 vccd1 _11298_/X sky130_fd_sc_hd__a21bo_1
XFILLER_79_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13037_ _13037_/A vssd1 vssd1 vccd1 vccd1 _13037_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_17914_ _18960_/CLK _17914_/D vssd1 vssd1 vccd1 vccd1 _17914_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_152_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10249_ _12074_/A vssd1 vssd1 vccd1 vccd1 _10829_/A sky130_fd_sc_hd__inv_2
XFILLER_39_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18894_ _18899_/CLK _18894_/D vssd1 vssd1 vccd1 vccd1 _18894_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_230_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_227_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17845_ _19021_/CLK _17845_/D vssd1 vssd1 vccd1 vccd1 _17845_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_67_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17776_ _19034_/Q _12228_/Y _12178_/X vssd1 vssd1 vccd1 vccd1 _19034_/D sky130_fd_sc_hd__o21a_1
X_14988_ _15232_/A vssd1 vssd1 vccd1 vccd1 _15042_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_35_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_223_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16727_ _16727_/A vssd1 vssd1 vccd1 vccd1 _16773_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_47_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_223_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13939_ _13434_/A _13931_/X _13938_/X _12055_/A vssd1 vssd1 vccd1 vccd1 _14009_/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_62_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_222_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16658_ _16699_/A _16658_/B vssd1 vssd1 vccd1 vccd1 _16658_/Y sky130_fd_sc_hd__nand2_1
XFILLER_62_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_223_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_179_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15609_ _15677_/A vssd1 vssd1 vccd1 vccd1 _15748_/C sky130_fd_sc_hd__buf_2
XFILLER_222_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16589_ _16634_/A _16589_/B vssd1 vssd1 vccd1 vccd1 _16589_/Y sky130_fd_sc_hd__nand2_1
XFILLER_124_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09130_ _18833_/Q _18832_/Q _18831_/Q vssd1 vssd1 vccd1 vccd1 _09131_/D sky130_fd_sc_hd__or3_4
XFILLER_194_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18328_ _18346_/CLK _18328_/D vssd1 vssd1 vccd1 vccd1 _18328_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_198_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_187_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09061_ _17838_/Q vssd1 vssd1 vccd1 vccd1 _09072_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_18259_ _18266_/CLK _18259_/D vssd1 vssd1 vccd1 vccd1 _18259_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_131_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09963_ _09360_/A _09370_/A _09365_/C _09360_/B _10291_/A _09950_/X vssd1 vssd1 vccd1
+ vccd1 _09964_/B sky130_fd_sc_hd__mux4_1
XFILLER_89_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_65_wb_clk_i clkbuf_5_21_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18677_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_134_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09894_ _09915_/A _12130_/A vssd1 vssd1 vccd1 vccd1 _09965_/A sky130_fd_sc_hd__and2_2
XFILLER_100_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_217_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_214_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_225_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09328_ _18533_/Q _18532_/Q _18531_/Q vssd1 vssd1 vccd1 vccd1 _09332_/A sky130_fd_sc_hd__or3_4
XFILLER_178_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_159_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09259_ _18959_/Q _18958_/Q _18957_/Q vssd1 vssd1 vccd1 vccd1 _09260_/D sky130_fd_sc_hd__or3_4
XFILLER_194_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_182_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12270_ _12270_/A _12270_/B vssd1 vssd1 vccd1 vccd1 _12289_/A sky130_fd_sc_hd__or2_2
XFILLER_154_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11221_ _11243_/A vssd1 vssd1 vccd1 vccd1 _11221_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_135_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_218_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11152_ _13509_/A vssd1 vssd1 vccd1 vccd1 _11584_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_68_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10103_ _10317_/A _10103_/B vssd1 vssd1 vccd1 vccd1 _10103_/X sky130_fd_sc_hd__or2_1
XFILLER_150_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15960_ _16003_/A _15960_/B vssd1 vssd1 vccd1 vccd1 _15960_/Y sky130_fd_sc_hd__nand2_1
XTAP_5410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11083_ _11083_/A vssd1 vssd1 vccd1 vccd1 _17790_/D sky130_fd_sc_hd__clkbuf_1
XTAP_5421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_191_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10034_ _09186_/A _09181_/A _09181_/D _09176_/D _09703_/A _12059_/A vssd1 vssd1 vccd1
+ vccd1 _10034_/X sky130_fd_sc_hd__mux4_2
X_14911_ _14913_/B _14909_/X _14910_/Y _14902_/X vssd1 vssd1 vccd1 vccd1 _18316_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_23_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15891_ _15890_/B _15888_/X _15890_/Y _15881_/X vssd1 vssd1 vccd1 vccd1 _18551_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_4720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17630_ _17630_/A vssd1 vssd1 vccd1 vccd1 _18970_/D sky130_fd_sc_hd__clkbuf_1
XTAP_5498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14842_ _18336_/Q _18300_/Q _14848_/S vssd1 vssd1 vccd1 vccd1 _14842_/X sky130_fd_sc_hd__mux2_1
XTAP_4764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_217_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17561_ _17675_/A vssd1 vssd1 vccd1 vccd1 _17561_/X sky130_fd_sc_hd__buf_2
X_14773_ _14793_/A _15371_/B _14818_/C vssd1 vssd1 vccd1 vccd1 _14773_/X sky130_fd_sc_hd__or3_1
X_11985_ _11985_/A _11985_/B _11988_/A _11985_/D vssd1 vssd1 vccd1 vccd1 _12009_/C
+ sky130_fd_sc_hd__or4_1
XFILLER_95_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_217_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_205_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16512_ _17119_/A _17119_/B _16512_/C _15903_/C vssd1 vssd1 vccd1 vccd1 _16976_/B
+ sky130_fd_sc_hd__or4b_4
X_13724_ _13724_/A vssd1 vssd1 vccd1 vccd1 _13743_/A sky130_fd_sc_hd__buf_4
XFILLER_95_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10936_ _10932_/X _10935_/X _10936_/S vssd1 vssd1 vccd1 vccd1 _10936_/X sky130_fd_sc_hd__mux2_1
XFILLER_44_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17492_ _18972_/Q _18936_/Q _17495_/S vssd1 vssd1 vccd1 vccd1 _17492_/X sky130_fd_sc_hd__mux2_1
XFILLER_210_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_182_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_231_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_189_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19231_ _19231_/A _08939_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[31] sky130_fd_sc_hd__ebufn_8
XFILLER_44_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16443_ _16503_/A vssd1 vssd1 vccd1 vccd1 _16491_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_13655_ _18972_/Q _13585_/A _13566_/A _18966_/Q vssd1 vssd1 vccd1 vccd1 _13655_/X
+ sky130_fd_sc_hd__a22o_1
X_10867_ _10867_/A _10867_/B vssd1 vssd1 vccd1 vccd1 _10867_/X sky130_fd_sc_hd__or2_1
XFILLER_223_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19162_ _19162_/A _09060_/Y vssd1 vssd1 vccd1 vccd1 io_out[0] sky130_fd_sc_hd__ebufn_8
X_12606_ _12608_/A _12609_/B vssd1 vssd1 vccd1 vccd1 _12607_/A sky130_fd_sc_hd__or2_1
X_16374_ _16891_/A vssd1 vssd1 vccd1 vccd1 _16780_/A sky130_fd_sc_hd__buf_2
X_13586_ _13586_/A vssd1 vssd1 vccd1 vccd1 _13856_/A sky130_fd_sc_hd__buf_2
XPHY_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10798_ _10779_/X _10793_/X _10797_/X _10910_/D vssd1 vssd1 vccd1 vccd1 _10798_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_223_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18113_ _18126_/CLK _18113_/D vssd1 vssd1 vccd1 vccd1 _18113_/Q sky130_fd_sc_hd__dfxtp_1
X_15325_ _15375_/A _15325_/B vssd1 vssd1 vccd1 vccd1 _15325_/Y sky130_fd_sc_hd__nand2_1
X_12537_ _12533_/Y _12535_/Y _12537_/S vssd1 vssd1 vccd1 vccd1 _12538_/B sky130_fd_sc_hd__mux2_1
XFILLER_185_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18044_ _18044_/CLK _18044_/D vssd1 vssd1 vccd1 vccd1 _18044_/Q sky130_fd_sc_hd__dfxtp_1
X_15256_ _18438_/Q _18402_/Q _15267_/S vssd1 vssd1 vccd1 vccd1 _15256_/X sky130_fd_sc_hd__mux2_1
X_12468_ _12468_/A vssd1 vssd1 vccd1 vccd1 _17905_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_173_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11419_ _17881_/Q vssd1 vssd1 vccd1 vccd1 _11419_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_14207_ _10985_/X _09709_/X _14205_/X _10413_/X _14206_/Y vssd1 vssd1 vccd1 vccd1
+ _14207_/X sky130_fd_sc_hd__a221o_1
X_15187_ _15187_/A vssd1 vssd1 vccd1 vccd1 _15187_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_141_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12399_ _12399_/A vssd1 vssd1 vccd1 vccd1 _17896_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_126_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14138_ _18344_/Q _13507_/A _13582_/A _18350_/Q vssd1 vssd1 vccd1 vccd1 _14138_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_141_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14069_ _18812_/Q _13591_/X _13861_/X _18836_/Q vssd1 vssd1 vccd1 vccd1 _14069_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_141_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18946_ _18950_/CLK _18946_/D vssd1 vssd1 vccd1 vccd1 _18946_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_140_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18877_ _18914_/CLK _18877_/D vssd1 vssd1 vccd1 vccd1 _18877_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_66_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17828_ _18157_/CLK _17828_/D vssd1 vssd1 vccd1 vccd1 _17828_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_82_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_227_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17759_ _17759_/A vssd1 vssd1 vccd1 vccd1 _19022_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_82_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_183_wb_clk_i clkbuf_5_9_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _19021_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_35_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_222_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_112_wb_clk_i clkbuf_5_30_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18504_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_74_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09113_ _18737_/Q _18736_/Q _18735_/Q vssd1 vssd1 vccd1 vccd1 _10728_/A sky130_fd_sc_hd__or3_4
XFILLER_109_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09044_ _09046_/A vssd1 vssd1 vccd1 vccd1 _09044_/Y sky130_fd_sc_hd__inv_2
XFILLER_159_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_159_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_209_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_132_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_213_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09946_ _09402_/A _09392_/B _09397_/C _10877_/A _09945_/X _09905_/X vssd1 vssd1 vccd1
+ vccd1 _09946_/X sky130_fd_sc_hd__mux4_2
XFILLER_89_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_213_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_11 _09153_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09877_ _10181_/A _09896_/B vssd1 vssd1 vccd1 vccd1 _09907_/A sky130_fd_sc_hd__nand2_2
XINSDIODE2_22 _09214_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_33 _09924_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_213_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_44 _10555_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_55 _15840_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_66 _13508_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_77 _13906_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_88 _13630_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_99 _13846_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11770_ _11770_/A _11770_/B _11770_/C vssd1 vssd1 vccd1 vccd1 _11776_/B sky130_fd_sc_hd__and3_1
XFILLER_198_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_1333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10721_ _10721_/A vssd1 vssd1 vccd1 vccd1 _10763_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_53_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_198_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_224_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13440_ _11984_/B _13426_/B _13439_/Y vssd1 vssd1 vccd1 vccd1 _13456_/B sky130_fd_sc_hd__a21o_1
XFILLER_9_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10652_ _10805_/A vssd1 vssd1 vccd1 vccd1 _10689_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_13_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_220_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13371_ _13371_/A vssd1 vssd1 vccd1 vccd1 _18108_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_194_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10583_ _09344_/C _09344_/D _09354_/D _09349_/D _09688_/A _09995_/A vssd1 vssd1 vccd1
+ vccd1 _10583_/X sky130_fd_sc_hd__mux4_2
XFILLER_70_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15110_ _18402_/Q _18366_/Q _15121_/S vssd1 vssd1 vccd1 vccd1 _15110_/X sky130_fd_sc_hd__mux2_1
X_12322_ _12333_/C _12327_/C vssd1 vssd1 vccd1 vccd1 _12323_/C sky130_fd_sc_hd__nor2_1
X_16090_ _16096_/B _16087_/X _16089_/X _16074_/X vssd1 vssd1 vccd1 vccd1 _18597_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_186_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_177_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15041_ _18384_/Q _18348_/Q _15052_/S vssd1 vssd1 vccd1 vccd1 _15041_/X sky130_fd_sc_hd__mux2_1
XFILLER_6_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12253_ _12253_/A _12258_/C vssd1 vssd1 vccd1 vccd1 _12253_/Y sky130_fd_sc_hd__nor2_1
XFILLER_218_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11204_ _11201_/A _11205_/C _17813_/Q vssd1 vssd1 vccd1 vccd1 _11206_/B sky130_fd_sc_hd__a21o_1
XFILLER_108_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12184_ _14436_/A vssd1 vssd1 vccd1 vccd1 _12184_/X sky130_fd_sc_hd__clkbuf_2
X_18800_ _18811_/CLK _18800_/D vssd1 vssd1 vccd1 vccd1 _18800_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_122_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11135_ _11582_/A vssd1 vssd1 vccd1 vccd1 _11661_/A sky130_fd_sc_hd__buf_2
XFILLER_122_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_231_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16992_ _17015_/A _17425_/B _17028_/C vssd1 vssd1 vccd1 vccd1 _16992_/X sky130_fd_sc_hd__or3_1
XFILLER_95_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18731_ _18765_/CLK _18731_/D vssd1 vssd1 vccd1 vccd1 _18731_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_135_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15943_ _15942_/B _15941_/X _15942_/Y _15925_/X vssd1 vssd1 vccd1 vccd1 _18563_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_5240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11066_ _11942_/A vssd1 vssd1 vccd1 vccd1 _11970_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_110_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_231_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10017_ _10015_/X _10016_/X _10017_/S vssd1 vssd1 vccd1 vccd1 _10017_/X sky130_fd_sc_hd__mux2_1
XTAP_5284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18662_ _18662_/CLK _18662_/D vssd1 vssd1 vccd1 vccd1 _18662_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_7_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15874_ _15876_/B _15872_/X _15873_/Y _15861_/X vssd1 vssd1 vccd1 vccd1 _18547_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_4550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17613_ _17571_/X _17602_/Y _17603_/X _17605_/Y _18965_/Q vssd1 vssd1 vccd1 vccd1
+ _17614_/B sky130_fd_sc_hd__a32o_1
XTAP_4583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14825_ _18332_/Q _18296_/Q _14830_/S vssd1 vssd1 vccd1 vccd1 _14825_/X sky130_fd_sc_hd__mux2_1
XFILLER_91_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_218_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18593_ _18593_/CLK _18593_/D vssd1 vssd1 vccd1 vccd1 _18593_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_221_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_224_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17544_ _17544_/A _17544_/B vssd1 vssd1 vccd1 vccd1 _17544_/Y sky130_fd_sc_hd__nand2_1
XTAP_3893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14756_ _18315_/Q _18279_/Q _14756_/S vssd1 vssd1 vccd1 vccd1 _14756_/X sky130_fd_sc_hd__mux2_1
X_11968_ _12023_/A _11974_/B _11999_/B _11929_/X _11281_/A vssd1 vssd1 vccd1 vccd1
+ _11968_/X sky130_fd_sc_hd__o311a_1
XFILLER_189_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_220_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13707_ _18753_/Q _14124_/A _13706_/X _18735_/Q vssd1 vssd1 vccd1 vccd1 _13707_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_205_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10919_ _09349_/D _09344_/D _09354_/D _09344_/C _10484_/X _10231_/X vssd1 vssd1 vccd1
+ vccd1 _10920_/B sky130_fd_sc_hd__mux4_2
X_17475_ _17509_/A _17477_/B vssd1 vssd1 vccd1 vccd1 _17475_/Y sky130_fd_sc_hd__nand2_1
X_14687_ _14687_/A _15277_/A vssd1 vssd1 vccd1 vccd1 _14700_/B sky130_fd_sc_hd__nor2_1
X_11899_ _17791_/Q _11951_/B _11899_/C vssd1 vssd1 vccd1 vccd1 _11947_/B sky130_fd_sc_hd__or3_2
XFILLER_220_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_220_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19214_ _19214_/A _08966_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[14] sky130_fd_sc_hd__ebufn_8
X_16426_ _16447_/A _16429_/B vssd1 vssd1 vccd1 vccd1 _16426_/Y sky130_fd_sc_hd__nand2_1
XFILLER_177_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13638_ _18900_/Q _13586_/A _13588_/A _18891_/Q vssd1 vssd1 vccd1 vccd1 _13638_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_220_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19145_ _19145_/A _09048_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[15] sky130_fd_sc_hd__ebufn_8
X_16357_ _18696_/Q _18660_/Q _16363_/S vssd1 vssd1 vccd1 vccd1 _16357_/X sky130_fd_sc_hd__mux2_1
XFILLER_160_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13569_ _18684_/Q _13621_/A _13568_/X _18678_/Q vssd1 vssd1 vccd1 vccd1 _13569_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_146_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15308_ _15440_/A vssd1 vssd1 vccd1 vccd1 _15415_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_160_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16288_ _16431_/A vssd1 vssd1 vccd1 vccd1 _16880_/B sky130_fd_sc_hd__buf_4
XFILLER_146_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18027_ _18030_/CLK _18027_/D vssd1 vssd1 vccd1 vccd1 _18027_/Q sky130_fd_sc_hd__dfxtp_1
X_15239_ _15239_/A _15239_/B vssd1 vssd1 vccd1 vccd1 _15239_/Y sky130_fd_sc_hd__nand2_1
XFILLER_172_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09800_ _09800_/A _09800_/B vssd1 vssd1 vccd1 vccd1 _09800_/X sky130_fd_sc_hd__and2_1
XFILLER_101_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_228_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09731_ _18102_/Q _17980_/Q vssd1 vssd1 vccd1 vccd1 _09732_/B sky130_fd_sc_hd__xor2_2
X_18929_ _18936_/CLK _18929_/D vssd1 vssd1 vccd1 vccd1 _18929_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_132_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_1232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09662_ _13372_/A _09623_/B _09661_/X vssd1 vssd1 vccd1 vccd1 _12080_/S sky130_fd_sc_hd__a21oi_2
XFILLER_27_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_215_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09593_ _09593_/A _09593_/B _09593_/C vssd1 vssd1 vccd1 vccd1 _09722_/B sky130_fd_sc_hd__or3_1
XFILLER_131_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_224_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_224_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_223_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_170 _18926_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_208_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINSDIODE2_181 _08972_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_211_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XINSDIODE2_192 _09143_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_168_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_80_wb_clk_i clkbuf_5_23_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18607_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_164_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09027_ _09028_/A vssd1 vssd1 vccd1 vccd1 _09027_/Y sky130_fd_sc_hd__inv_2
XFILLER_151_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09929_ _12122_/A _12130_/A vssd1 vssd1 vccd1 vccd1 _09930_/A sky130_fd_sc_hd__nor2_2
XFILLER_120_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_218_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12940_ _12940_/A vssd1 vssd1 vccd1 vccd1 _13049_/A sky130_fd_sc_hd__buf_2
XTAP_3101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_213_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12871_ _12871_/A _12871_/B vssd1 vssd1 vccd1 vccd1 _12877_/C sky130_fd_sc_hd__nor2_1
XFILLER_73_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14610_ _14915_/A vssd1 vssd1 vccd1 vccd1 _17471_/A sky130_fd_sc_hd__buf_8
XTAP_3178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11822_ _17556_/A vssd1 vssd1 vccd1 vccd1 _11822_/X sky130_fd_sc_hd__buf_6
XTAP_2444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15590_ _18514_/Q _18478_/Q _15604_/S vssd1 vssd1 vccd1 vccd1 _15590_/X sky130_fd_sc_hd__mux2_1
XTAP_1710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11753_ _11753_/A _11760_/B vssd1 vssd1 vccd1 vccd1 _11753_/X sky130_fd_sc_hd__or2_1
X_14541_ _18184_/Q vssd1 vssd1 vccd1 vccd1 _15957_/A sky130_fd_sc_hd__inv_2
XTAP_2488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10704_ _10867_/A _10703_/X _10679_/A vssd1 vssd1 vccd1 vccd1 _10704_/X sky130_fd_sc_hd__a21o_1
XFILLER_183_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17260_ _17304_/A vssd1 vssd1 vccd1 vccd1 _17260_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_109_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11684_ _19033_/Q vssd1 vssd1 vccd1 vccd1 _11696_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_14472_ _14472_/A vssd1 vssd1 vccd1 vccd1 _18210_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16211_ _18661_/Q _18625_/Q _16215_/S vssd1 vssd1 vccd1 vccd1 _16211_/X sky130_fd_sc_hd__mux2_1
XFILLER_139_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13423_ _13648_/A _13649_/B vssd1 vssd1 vccd1 vccd1 _13710_/C sky130_fd_sc_hd__or2_4
X_10635_ _12966_/A _10650_/B _12074_/A vssd1 vssd1 vccd1 vccd1 _10654_/A sky130_fd_sc_hd__a21oi_2
X_17191_ _17480_/A _17202_/B vssd1 vssd1 vccd1 vccd1 _17200_/B sky130_fd_sc_hd__nor2_2
XFILLER_128_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_1366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16142_ _16212_/A vssd1 vssd1 vccd1 vccd1 _16199_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_167_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13354_ _13346_/X _13353_/Y _11023_/X vssd1 vssd1 vccd1 vccd1 _18104_/D sky130_fd_sc_hd__a21boi_1
X_10566_ _09304_/A _09294_/B _09299_/C _09304_/C _10089_/S _10036_/X vssd1 vssd1 vccd1
+ vccd1 _10566_/X sky130_fd_sc_hd__mux4_2
XFILLER_220_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_194_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_182_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12305_ _11218_/X _11385_/B _12304_/Y _12313_/B _11323_/B vssd1 vssd1 vccd1 vccd1
+ _17876_/D sky130_fd_sc_hd__a32o_1
XFILLER_155_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16073_ _16115_/A _16678_/B _16115_/C vssd1 vssd1 vccd1 vccd1 _16073_/X sky130_fd_sc_hd__or3_1
X_13285_ _18025_/Q _18024_/Q _18027_/Q _18026_/Q vssd1 vssd1 vccd1 vccd1 _13286_/D
+ sky130_fd_sc_hd__or4_1
XFILLER_170_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10497_ _09098_/A _09103_/D _10550_/S vssd1 vssd1 vccd1 vccd1 _10497_/X sky130_fd_sc_hd__mux2_1
XFILLER_120_1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15024_ _18380_/Q _18344_/Q _15033_/S vssd1 vssd1 vccd1 vccd1 _15024_/X sky130_fd_sc_hd__mux2_1
XFILLER_154_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12236_ _17859_/Q _11603_/A _12223_/X vssd1 vssd1 vccd1 vccd1 _12246_/A sky130_fd_sc_hd__o21ai_1
XFILLER_114_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_170_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12167_ _12160_/Y _12166_/X _12163_/X vssd1 vssd1 vccd1 vccd1 _17844_/D sky130_fd_sc_hd__o21a_1
XFILLER_123_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11118_ _11788_/A vssd1 vssd1 vccd1 vccd1 _11735_/A sky130_fd_sc_hd__clkbuf_2
X_12098_ _14330_/A _13710_/A vssd1 vssd1 vccd1 vccd1 _12104_/C sky130_fd_sc_hd__xnor2_1
X_16975_ _16975_/A vssd1 vssd1 vccd1 vccd1 _16975_/X sky130_fd_sc_hd__buf_2
XFILLER_96_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18714_ _18722_/CLK _18714_/D vssd1 vssd1 vccd1 vccd1 _18714_/Q sky130_fd_sc_hd__dfxtp_1
X_15926_ _15928_/B _15923_/X _15924_/Y _15925_/X vssd1 vssd1 vccd1 vccd1 _18559_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_5070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11049_ _11042_/X _09802_/B _11026_/X _11045_/X _13383_/A vssd1 vssd1 vccd1 vccd1
+ _17784_/D sky130_fd_sc_hd__o2111a_1
XFILLER_77_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_225_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18645_ _18683_/CLK _18645_/D vssd1 vssd1 vccd1 vccd1 _18645_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_76_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15857_ _15857_/A _16007_/B _15870_/C vssd1 vssd1 vccd1 vccd1 _15857_/X sky130_fd_sc_hd__or3_1
XTAP_4380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14808_ _14814_/B _14805_/X _14807_/X _14799_/X vssd1 vssd1 vccd1 vccd1 _18291_/D
+ sky130_fd_sc_hd__o211a_1
X_18576_ _18577_/CLK _18576_/D vssd1 vssd1 vccd1 vccd1 _18576_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_92_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15788_ _15799_/A _15935_/B _15811_/C vssd1 vssd1 vccd1 vccd1 _15788_/X sky130_fd_sc_hd__or3_1
XTAP_3690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_229_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17527_ _18981_/Q _18945_/Q _17533_/S vssd1 vssd1 vccd1 vccd1 _17527_/X sky130_fd_sc_hd__mux2_1
XFILLER_221_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14739_ _14742_/B _14736_/X _14737_/Y _14738_/X vssd1 vssd1 vccd1 vccd1 _18274_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_33_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17458_ _17458_/A _17491_/B vssd1 vssd1 vccd1 vccd1 _17469_/B sky130_fd_sc_hd__nor2_2
XFILLER_178_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16409_ _16701_/A _16452_/B vssd1 vssd1 vccd1 vccd1 _16417_/B sky130_fd_sc_hd__nor2_1
XFILLER_193_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_220_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_203_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17389_ _17395_/B _17386_/X _17388_/X _17380_/X vssd1 vssd1 vccd1 vccd1 _18909_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_9_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_1321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_206_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_214_1362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_228_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09714_ _18254_/Q _18253_/Q _18252_/Q vssd1 vssd1 vccd1 vccd1 _09714_/X sky130_fd_sc_hd__or3_4
XFILLER_142_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_228_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_216_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09645_ _09645_/A _09645_/B vssd1 vssd1 vccd1 vccd1 _09647_/B sky130_fd_sc_hd__xnor2_1
XFILLER_215_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_222_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09576_ _09600_/A _09576_/B vssd1 vssd1 vccd1 vccd1 _09585_/B sky130_fd_sc_hd__nor2_1
XTAP_1017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_231_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_224_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_2_0_0_wb_clk_i clkbuf_2_1_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_2_0_1_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_23_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_204_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10420_ _09209_/B _09219_/C _09219_/D _09214_/A _10236_/A _10413_/X vssd1 vssd1 vccd1
+ vccd1 _10420_/X sky130_fd_sc_hd__mux4_2
XFILLER_17_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_183_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10351_ _09114_/C _09950_/X _10350_/X _09969_/A vssd1 vssd1 vccd1 vccd1 _10351_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_136_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_1216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_178_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_191_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13070_ _14421_/A _13070_/B vssd1 vssd1 vccd1 vccd1 _13071_/A sky130_fd_sc_hd__or2_1
X_10282_ _09170_/B _09160_/B _10286_/S vssd1 vssd1 vccd1 vccd1 _10282_/X sky130_fd_sc_hd__mux2_1
XFILLER_133_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12021_ _12021_/A _12021_/B vssd1 vssd1 vccd1 vccd1 _12042_/A sky130_fd_sc_hd__nor2_8
XFILLER_120_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_215_wb_clk_i clkbuf_5_8_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17888_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_104_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16760_ _16760_/A vssd1 vssd1 vccd1 vccd1 _16760_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_24_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13972_ _18289_/Q _13848_/A _13654_/X _18280_/Q _13971_/X vssd1 vssd1 vccd1 vccd1
+ _13972_/X sky130_fd_sc_hd__a221o_1
XFILLER_24_1176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15711_ _18543_/Q _18507_/Q _15714_/S vssd1 vssd1 vccd1 vccd1 _15711_/X sky130_fd_sc_hd__mux2_1
XFILLER_207_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12923_ _18000_/Q _12770_/Y _18036_/Q _12919_/X _12983_/A vssd1 vssd1 vccd1 vccd1
+ _12923_/Y sky130_fd_sc_hd__a41oi_1
XFILLER_46_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16691_ _16808_/A vssd1 vssd1 vccd1 vccd1 _16736_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_207_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18430_ _18434_/CLK _18430_/D vssd1 vssd1 vccd1 vccd1 _18430_/Q sky130_fd_sc_hd__dfxtp_4
X_15642_ _18526_/Q _18490_/Q _15642_/S vssd1 vssd1 vccd1 vccd1 _15642_/X sky130_fd_sc_hd__mux2_1
XFILLER_62_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12854_ _12874_/A vssd1 vssd1 vccd1 vccd1 _12854_/X sky130_fd_sc_hd__buf_2
XTAP_2241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_222_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18361_ _18393_/CLK _18361_/D vssd1 vssd1 vccd1 vccd1 _18361_/Q sky130_fd_sc_hd__dfxtp_4
X_11805_ _11070_/X _11312_/B _11964_/A vssd1 vssd1 vccd1 vccd1 _11808_/C sky130_fd_sc_hd__o21a_1
XTAP_2274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15573_ _18510_/Q _18474_/Q _15586_/S vssd1 vssd1 vccd1 vccd1 _15573_/X sky130_fd_sc_hd__mux2_1
XFILLER_15_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12785_ _17942_/Q _12776_/X _12784_/X _12318_/X vssd1 vssd1 vccd1 vccd1 _17942_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_61_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17312_ _17314_/B _17310_/X _17311_/Y _17304_/X vssd1 vssd1 vccd1 vccd1 _18889_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_15_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14524_ _18180_/Q _18179_/Q _18181_/Q vssd1 vssd1 vccd1 vccd1 _14704_/C sky130_fd_sc_hd__nand3b_2
XFILLER_230_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18292_ _18312_/CLK _18292_/D vssd1 vssd1 vccd1 vccd1 _18292_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_15_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11736_ _17913_/Q vssd1 vssd1 vccd1 vccd1 _11767_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_202_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17243_ _17526_/A _17254_/B vssd1 vssd1 vccd1 vccd1 _17252_/B sky130_fd_sc_hd__nor2_1
X_14455_ _17766_/A _14455_/B vssd1 vssd1 vccd1 vccd1 _18204_/D sky130_fd_sc_hd__nor2_1
X_11667_ _12251_/A _11671_/B _11651_/A vssd1 vssd1 vccd1 vccd1 _11668_/B sky130_fd_sc_hd__o21a_1
XFILLER_179_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13406_ _13406_/A vssd1 vssd1 vccd1 vccd1 _18128_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_127_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10618_ _10618_/A vssd1 vssd1 vccd1 vccd1 _10619_/A sky130_fd_sc_hd__inv_2
X_17174_ _17180_/B _17172_/X _17173_/X _17161_/X vssd1 vssd1 vccd1 vccd1 _18855_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_128_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11598_ _11868_/B _11598_/B vssd1 vssd1 vccd1 vccd1 _11850_/A sky130_fd_sc_hd__nand2_1
X_14386_ _14386_/A _14386_/B vssd1 vssd1 vccd1 vccd1 _14386_/Y sky130_fd_sc_hd__nor2_2
XFILLER_155_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16125_ _16287_/A _16208_/C vssd1 vssd1 vccd1 vccd1 _16132_/B sky130_fd_sc_hd__nor2_2
X_10549_ _10549_/A _10549_/B vssd1 vssd1 vccd1 vccd1 _10549_/X sky130_fd_sc_hd__or2_1
XFILLER_115_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13337_ _13337_/A vssd1 vssd1 vccd1 vccd1 _13337_/X sky130_fd_sc_hd__buf_2
XFILLER_182_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16056_ _16193_/A vssd1 vssd1 vccd1 vccd1 _16115_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_192_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13268_ _13467_/A input4/X vssd1 vssd1 vccd1 vccd1 _18087_/D sky130_fd_sc_hd__nor2_1
XFILLER_68_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15007_ _15247_/A vssd1 vssd1 vccd1 vccd1 _15058_/A sky130_fd_sc_hd__buf_2
X_12219_ _13037_/A vssd1 vssd1 vccd1 vccd1 _12219_/X sky130_fd_sc_hd__buf_6
XFILLER_69_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13199_ _13199_/A vssd1 vssd1 vccd1 vccd1 _13208_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_96_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16958_ _16957_/B _16956_/X _16957_/Y _16940_/X vssd1 vssd1 vccd1 vccd1 _18803_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_49_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15909_ _15921_/A _15909_/B _15964_/C vssd1 vssd1 vccd1 vccd1 _15909_/X sky130_fd_sc_hd__or3_1
X_16889_ _16889_/A vssd1 vssd1 vccd1 vccd1 _17483_/B sky130_fd_sc_hd__buf_6
XFILLER_225_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09430_ _09188_/X _09428_/X _09430_/C _09430_/D vssd1 vssd1 vccd1 vccd1 _09470_/A
+ sky130_fd_sc_hd__and4bb_1
X_18628_ _18658_/CLK _18628_/D vssd1 vssd1 vccd1 vccd1 _18628_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_25_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_225_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_213_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09361_ _18272_/Q _18271_/Q _18270_/Q vssd1 vssd1 vccd1 vccd1 _09365_/A sky130_fd_sc_hd__or3_2
X_18559_ _18572_/CLK _18559_/D vssd1 vssd1 vccd1 vccd1 _18559_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_24_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_19_wb_clk_i clkbuf_5_5_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18907_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_09292_ _18506_/Q _18505_/Q _18504_/Q vssd1 vssd1 vccd1 vccd1 _09294_/C sky130_fd_sc_hd__or3_4
XFILLER_75_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_1364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_203_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_133_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_217_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_1293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_228_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_216_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_216_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09628_ _13372_/A _09631_/B _09627_/X vssd1 vssd1 vccd1 vccd1 _09665_/B sky130_fd_sc_hd__a21oi_2
XFILLER_189_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09559_ _10044_/A vssd1 vssd1 vccd1 vccd1 _10895_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_197_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_1272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_197_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12570_ _17923_/Q _12570_/B vssd1 vssd1 vccd1 vccd1 _12570_/Y sky130_fd_sc_hd__nor2_1
XFILLER_52_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_212_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11521_ _17871_/Q _17870_/Q vssd1 vssd1 vccd1 vccd1 _12285_/C sky130_fd_sc_hd__nand2_1
XFILLER_196_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11452_ _11452_/A _11788_/B vssd1 vssd1 vccd1 vccd1 _13429_/A sky130_fd_sc_hd__or2_4
X_14240_ _14260_/A _14240_/B vssd1 vssd1 vccd1 vccd1 _14240_/Y sky130_fd_sc_hd__nand2_1
XFILLER_172_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_184_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10403_ _10403_/A _10403_/B _10366_/B vssd1 vssd1 vccd1 vccd1 _10403_/X sky130_fd_sc_hd__or3b_1
X_14171_ _18596_/Q _14019_/X _14030_/X _18620_/Q vssd1 vssd1 vccd1 vccd1 _14171_/X
+ sky130_fd_sc_hd__a22o_1
X_11383_ _12299_/B _11828_/A _11378_/Y _11379_/X _11619_/A vssd1 vssd1 vccd1 vccd1
+ _11384_/A sky130_fd_sc_hd__o32a_1
XFILLER_109_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13122_ _13122_/A vssd1 vssd1 vccd1 vccd1 _18020_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_3_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10334_ _09889_/X _10330_/X _10333_/X _09981_/A vssd1 vssd1 vccd1 vccd1 _10334_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_194_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_180_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13053_ _13085_/A _18003_/Q _18005_/Q vssd1 vssd1 vccd1 vccd1 _13055_/B sky130_fd_sc_hd__a21boi_1
X_17930_ _17933_/CLK _17930_/D vssd1 vssd1 vccd1 vccd1 _17930_/Q sky130_fd_sc_hd__dfxtp_1
X_10265_ _10923_/S _10245_/X _10513_/A vssd1 vssd1 vccd1 vccd1 _10265_/X sky130_fd_sc_hd__a21bo_1
XFILLER_127_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12004_ _12025_/A _12026_/C vssd1 vssd1 vccd1 vccd1 _12004_/Y sky130_fd_sc_hd__nand2_1
XFILLER_121_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17861_ _17861_/CLK _17861_/D vssd1 vssd1 vccd1 vccd1 _17861_/Q sky130_fd_sc_hd__dfxtp_1
X_10196_ _13353_/A _10204_/B _10195_/X vssd1 vssd1 vccd1 vccd1 _10197_/B sky130_fd_sc_hd__a21oi_2
X_16812_ _18771_/Q _16815_/B _16811_/X _16800_/X vssd1 vssd1 vccd1 vccd1 _18771_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_93_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17792_ _17793_/CLK _17792_/D vssd1 vssd1 vccd1 vccd1 _17792_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_226_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16743_ _16755_/A _16743_/B vssd1 vssd1 vccd1 vccd1 _16743_/Y sky130_fd_sc_hd__nand2_1
XFILLER_115_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13955_ _12027_/C _13947_/X _13954_/X _12028_/A vssd1 vssd1 vccd1 vccd1 _14009_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_74_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12906_ _12908_/B _12915_/B _12906_/C vssd1 vssd1 vccd1 vccd1 _12907_/A sky130_fd_sc_hd__and3b_1
XFILLER_98_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16674_ _18137_/Q _17278_/B vssd1 vssd1 vccd1 vccd1 _16787_/A sky130_fd_sc_hd__nand2_1
XFILLER_19_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13886_ _18955_/Q _13642_/A _13513_/A _18961_/Q vssd1 vssd1 vccd1 vccd1 _13886_/X
+ sky130_fd_sc_hd__a22o_1
X_18413_ _18432_/CLK _18413_/D vssd1 vssd1 vccd1 vccd1 _18413_/Q sky130_fd_sc_hd__dfxtp_2
X_15625_ _16566_/A vssd1 vssd1 vccd1 vccd1 _15869_/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12837_ _12847_/A vssd1 vssd1 vccd1 vccd1 _12874_/A sky130_fd_sc_hd__clkbuf_2
XTAP_2071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18344_ _18346_/CLK _18344_/D vssd1 vssd1 vccd1 vccd1 _18344_/Q sky130_fd_sc_hd__dfxtp_2
X_15556_ _15558_/B _15553_/X _15554_/Y _15555_/X vssd1 vssd1 vccd1 vccd1 _18469_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_163_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12768_ _12987_/A _18993_/Q vssd1 vssd1 vccd1 vccd1 _12924_/B sky130_fd_sc_hd__or2_1
XTAP_1381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14507_ _14507_/A _14507_/B vssd1 vssd1 vccd1 vccd1 _14513_/B sky130_fd_sc_hd__or2_1
XFILLER_72_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_230_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18275_ _18275_/CLK _18275_/D vssd1 vssd1 vccd1 vccd1 _18275_/Q sky130_fd_sc_hd__dfxtp_1
X_11719_ _11720_/A _11719_/B vssd1 vssd1 vccd1 vccd1 _11742_/B sky130_fd_sc_hd__and2_1
X_15487_ _15511_/A _15487_/B vssd1 vssd1 vccd1 vccd1 _15487_/Y sky130_fd_sc_hd__nand2_1
XFILLER_148_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12699_ _17938_/Q vssd1 vssd1 vccd1 vccd1 _12699_/Y sky130_fd_sc_hd__inv_2
X_17226_ _17226_/A vssd1 vssd1 vccd1 vccd1 _17244_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_30_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14438_ _18200_/Q vssd1 vssd1 vccd1 vccd1 _14438_/Y sky130_fd_sc_hd__inv_2
XFILLER_175_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_128_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17157_ _17156_/B _17155_/X _17156_/Y _17140_/X vssd1 vssd1 vccd1 vccd1 _18851_/D
+ sky130_fd_sc_hd__o211a_1
X_14369_ _18186_/Q _18185_/Q _14381_/A vssd1 vssd1 vccd1 vccd1 _14375_/B sky130_fd_sc_hd__or3_1
XFILLER_157_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16108_ _18638_/Q _18602_/Q _16113_/S vssd1 vssd1 vccd1 vccd1 _16108_/X sky130_fd_sc_hd__mux2_1
XFILLER_192_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_137_wb_clk_i clkbuf_5_27_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18367_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_155_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17088_ _17088_/A _17091_/B vssd1 vssd1 vccd1 vccd1 _17088_/Y sky130_fd_sc_hd__nand2_1
X_19124__95 vssd1 vssd1 vccd1 vccd1 _19124__95/HI _19232_/A sky130_fd_sc_hd__conb_1
XFILLER_115_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16039_ _16064_/A _16039_/B vssd1 vssd1 vccd1 vccd1 _16039_/Y sky130_fd_sc_hd__nand2_1
X_08930_ _11018_/A vssd1 vssd1 vccd1 vccd1 _08935_/A sky130_fd_sc_hd__buf_12
XFILLER_83_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_229_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_1354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_226_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09413_ _09413_/A _10956_/A _09413_/C _09413_/D vssd1 vssd1 vccd1 vccd1 _09419_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_25_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_197_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_213_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09344_ _09344_/A _09344_/B _09344_/C _09344_/D vssd1 vssd1 vccd1 vccd1 _09355_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_90_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09275_ _18854_/Q _18853_/Q _18852_/Q vssd1 vssd1 vccd1 vccd1 _09277_/C sky130_fd_sc_hd__or3_2
XFILLER_32_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10050_ _09170_/A _09165_/D _09160_/D _09170_/C _09682_/A _09986_/A vssd1 vssd1 vccd1
+ vccd1 _10050_/X sky130_fd_sc_hd__mux4_1
XFILLER_88_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_229_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_217_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_216_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13740_ _18324_/Q _13585_/A _13739_/X _18315_/Q vssd1 vssd1 vccd1 vccd1 _13740_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_16_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10952_ _10962_/A _10952_/B vssd1 vssd1 vccd1 vccd1 _10952_/X sky130_fd_sc_hd__or2_1
XFILLER_43_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_1326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13671_ _13724_/A vssd1 vssd1 vccd1 vccd1 _13766_/A sky130_fd_sc_hd__buf_6
X_10883_ _10883_/A _10883_/B vssd1 vssd1 vccd1 vccd1 _10883_/X sky130_fd_sc_hd__or2_1
X_15410_ _15423_/A _16007_/B _15423_/C vssd1 vssd1 vccd1 vccd1 _15410_/X sky130_fd_sc_hd__or3_1
XFILLER_189_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12622_ _12629_/A _12569_/X _12619_/X _12620_/Y _12621_/X vssd1 vssd1 vccd1 vccd1
+ _17926_/D sky130_fd_sc_hd__a221o_1
XPHY_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16390_ _16392_/B _16388_/X _16389_/Y _16376_/X vssd1 vssd1 vccd1 vccd1 _18667_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_19_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_231_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_223_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15341_ _15339_/B _15338_/X _15339_/Y _15340_/X vssd1 vssd1 vccd1 vccd1 _18419_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_129_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12553_ _12588_/B _17919_/Q vssd1 vssd1 vccd1 vccd1 _12554_/B sky130_fd_sc_hd__and2_1
XFILLER_169_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_223_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_184_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11504_ _11412_/A _11617_/C _11594_/A _11412_/C vssd1 vssd1 vccd1 vccd1 _11504_/X
+ sky130_fd_sc_hd__o31a_1
X_18060_ _18072_/CLK _18060_/D vssd1 vssd1 vccd1 vccd1 _18060_/Q sky130_fd_sc_hd__dfxtp_1
X_15272_ _15301_/A _15275_/B vssd1 vssd1 vccd1 vccd1 _15272_/Y sky130_fd_sc_hd__nand2_1
XFILLER_106_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12484_ _12484_/A _12484_/B vssd1 vssd1 vccd1 vccd1 _12484_/X sky130_fd_sc_hd__or2_1
XFILLER_8_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_184_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17011_ _17010_/B _17009_/X _17010_/Y _16999_/X vssd1 vssd1 vccd1 vccd1 _18815_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_8_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14223_ _18206_/Q vssd1 vssd1 vccd1 vccd1 _14279_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_171_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11435_ _12316_/B _11377_/A _11432_/Y _11434_/X _11828_/B vssd1 vssd1 vccd1 vccd1
+ _11436_/A sky130_fd_sc_hd__o32a_1
XFILLER_7_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_230_wb_clk_i clkbuf_5_0_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17911_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_171_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14154_ _18758_/Q _13856_/X _13493_/X _18749_/Q _14153_/X vssd1 vssd1 vccd1 vccd1
+ _14154_/X sky130_fd_sc_hd__a221o_1
XFILLER_152_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11366_ _11366_/A _11843_/B vssd1 vssd1 vccd1 vccd1 _11577_/B sky130_fd_sc_hd__or2_1
XFILLER_98_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_217_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_152_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13105_ _13107_/A _18014_/Q vssd1 vssd1 vccd1 vccd1 _13106_/A sky130_fd_sc_hd__and2_1
X_10317_ _10317_/A _10599_/S vssd1 vssd1 vccd1 vccd1 _10317_/X sky130_fd_sc_hd__or2_1
XFILLER_153_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14085_ _18452_/Q _13508_/X _13842_/X _18458_/Q _14084_/X vssd1 vssd1 vccd1 vccd1
+ _14085_/X sky130_fd_sc_hd__a221o_1
X_11297_ _11313_/B _11297_/B _11297_/C vssd1 vssd1 vccd1 vccd1 _11297_/Y sky130_fd_sc_hd__nand3b_4
X_18962_ _18972_/CLK _18962_/D vssd1 vssd1 vccd1 vccd1 _18962_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_65_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13036_ _17991_/Q _13036_/B vssd1 vssd1 vccd1 vccd1 _13036_/X sky130_fd_sc_hd__or2_1
X_17913_ _18960_/CLK _17913_/D vssd1 vssd1 vccd1 vccd1 _17913_/Q sky130_fd_sc_hd__dfxtp_2
X_10248_ _17976_/Q vssd1 vssd1 vccd1 vccd1 _12074_/A sky130_fd_sc_hd__buf_2
XFILLER_117_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18893_ _18893_/CLK _18893_/D vssd1 vssd1 vccd1 vccd1 _18893_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_6_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_230_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17844_ _19019_/CLK _17844_/D vssd1 vssd1 vccd1 vccd1 _17844_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_227_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10179_ _10179_/A _10179_/B vssd1 vssd1 vccd1 vccd1 _12047_/A sky130_fd_sc_hd__xnor2_4
XFILLER_152_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17775_ _11696_/C _12205_/X _12178_/X vssd1 vssd1 vccd1 vccd1 _19033_/D sky130_fd_sc_hd__o21a_1
XFILLER_226_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14987_ _17575_/A vssd1 vssd1 vccd1 vccd1 _15232_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_19_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16726_ _17037_/A _16796_/C vssd1 vssd1 vccd1 vccd1 _16732_/B sky130_fd_sc_hd__nor2_2
X_13938_ _18337_/Q _13730_/X _13732_/X _18328_/Q _13937_/X vssd1 vssd1 vccd1 vccd1
+ _13938_/X sky130_fd_sc_hd__a221o_2
XFILLER_34_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_222_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_223_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_228_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_223_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16657_ _18770_/Q _18734_/Q _16657_/S vssd1 vssd1 vccd1 vccd1 _16657_/X sky130_fd_sc_hd__mux2_1
X_13869_ _13869_/A vssd1 vssd1 vccd1 vccd1 _14019_/A sky130_fd_sc_hd__buf_6
XFILLER_90_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_222_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15608_ _15757_/A _17410_/A vssd1 vssd1 vccd1 vccd1 _15677_/A sky130_fd_sc_hd__or2_1
XFILLER_179_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16588_ _16832_/A vssd1 vssd1 vccd1 vccd1 _16634_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_222_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18327_ _18346_/CLK _18327_/D vssd1 vssd1 vccd1 vccd1 _18327_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_124_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15539_ _18501_/Q _18465_/Q _15545_/S vssd1 vssd1 vccd1 vccd1 _15539_/X sky130_fd_sc_hd__mux2_1
XFILLER_188_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_1292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_202_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_176_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09060_ _11018_/A vssd1 vssd1 vccd1 vccd1 _09060_/Y sky130_fd_sc_hd__inv_2
XFILLER_175_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18258_ _18266_/CLK _18258_/D vssd1 vssd1 vccd1 vccd1 _18258_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_163_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17209_ _18901_/Q _18865_/Q _17221_/S vssd1 vssd1 vccd1 vccd1 _17209_/X sky130_fd_sc_hd__mux2_1
XFILLER_175_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18189_ _18191_/CLK _18189_/D vssd1 vssd1 vccd1 vccd1 _18189_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_190_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09962_ _09962_/A vssd1 vssd1 vccd1 vccd1 _10291_/A sky130_fd_sc_hd__buf_8
XFILLER_98_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09893_ _09920_/B vssd1 vssd1 vccd1 vccd1 _12130_/A sky130_fd_sc_hd__clkbuf_4
XTAP_951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_214_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_226_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_34_wb_clk_i clkbuf_5_18_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18244_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_26_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_225_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_167_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09327_ _09327_/A _09327_/B _09327_/C _09327_/D vssd1 vssd1 vccd1 vccd1 _09338_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_142_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_159_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09258_ _18953_/Q _18952_/Q _18951_/Q vssd1 vssd1 vccd1 vccd1 _10317_/A sky130_fd_sc_hd__or3_2
XFILLER_194_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_182_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09189_ _18560_/Q _18559_/Q _18558_/Q vssd1 vssd1 vccd1 vccd1 _09193_/A sky130_fd_sc_hd__or3_4
XFILLER_166_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11220_ _11224_/C _11220_/B vssd1 vssd1 vccd1 vccd1 _17816_/D sky130_fd_sc_hd__nor2_1
XFILLER_175_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_190_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11151_ _17803_/Q vssd1 vssd1 vccd1 vccd1 _13509_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_108_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10102_ _09270_/B _09260_/D _10102_/S vssd1 vssd1 vccd1 vccd1 _10102_/X sky130_fd_sc_hd__mux2_1
XFILLER_161_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11082_ _11334_/A _11232_/B _11091_/S vssd1 vssd1 vccd1 vccd1 _11083_/A sky130_fd_sc_hd__mux2_1
XFILLER_122_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_216_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14910_ _14932_/A _14913_/B vssd1 vssd1 vccd1 vccd1 _14910_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10033_ _10033_/A vssd1 vssd1 vccd1 vccd1 _14317_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_88_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_216_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15890_ _15942_/A _15890_/B vssd1 vssd1 vccd1 vccd1 _15890_/Y sky130_fd_sc_hd__nand2_1
XTAP_4710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14841_ _15277_/A _14841_/B vssd1 vssd1 vccd1 vccd1 _14849_/B sky130_fd_sc_hd__nor2_2
XFILLER_114_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17560_ _17602_/A _17635_/A vssd1 vssd1 vccd1 vccd1 _17560_/Y sky130_fd_sc_hd__nor2_2
XFILLER_84_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14772_ _14772_/A vssd1 vssd1 vccd1 vccd1 _14818_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_223_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_217_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11984_ _12023_/A _11984_/B _11984_/C vssd1 vssd1 vccd1 vccd1 _11985_/D sky130_fd_sc_hd__and3b_1
XFILLER_112_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16511_ _16510_/B _16509_/X _16510_/Y _16496_/X vssd1 vssd1 vccd1 vccd1 _18698_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_186_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13723_ _13741_/A vssd1 vssd1 vccd1 vccd1 _13723_/X sky130_fd_sc_hd__buf_6
X_10935_ _10933_/X _10934_/X _10935_/S vssd1 vssd1 vccd1 vccd1 _10935_/X sky130_fd_sc_hd__mux2_2
X_17491_ _17491_/A _17491_/B vssd1 vssd1 vccd1 vccd1 _17501_/B sky130_fd_sc_hd__nor2_2
XFILLER_17_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19230_ _19230_/A _08944_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[30] sky130_fd_sc_hd__ebufn_8
XFILLER_44_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16442_ _18717_/Q _18681_/Q _16449_/S vssd1 vssd1 vccd1 vccd1 _16442_/X sky130_fd_sc_hd__mux2_1
XFILLER_204_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_231_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13654_ _13654_/A vssd1 vssd1 vccd1 vccd1 _13654_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_31_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10866_ _09712_/X _09713_/X _09714_/X _09715_/X _10856_/S _14206_/A vssd1 vssd1 vccd1
+ vccd1 _10867_/B sky130_fd_sc_hd__mux4_2
XFILLER_143_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19161_ _19161_/A _09025_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[31] sky130_fd_sc_hd__ebufn_8
XPHY_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12605_ _17928_/Q vssd1 vssd1 vccd1 vccd1 _12608_/A sky130_fd_sc_hd__inv_2
XFILLER_231_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_223_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16373_ _16389_/A _16378_/B vssd1 vssd1 vccd1 vccd1 _16373_/Y sky130_fd_sc_hd__nand2_1
XPHY_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13585_ _13585_/A vssd1 vssd1 vccd1 vccd1 _13586_/A sky130_fd_sc_hd__buf_4
XPHY_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10797_ _10702_/A _10794_/X _10796_/X _10801_/S vssd1 vssd1 vccd1 vccd1 _10797_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_34_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18112_ _18125_/CLK _18112_/D vssd1 vssd1 vccd1 vccd1 _18112_/Q sky130_fd_sc_hd__dfxtp_1
X_15324_ _15582_/A vssd1 vssd1 vccd1 vccd1 _15375_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_169_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_184_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12536_ _12591_/A vssd1 vssd1 vccd1 vccd1 _12537_/S sky130_fd_sc_hd__buf_2
XFILLER_173_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18043_ _18094_/CLK _18043_/D vssd1 vssd1 vccd1 vccd1 _18043_/Q sky130_fd_sc_hd__dfxtp_1
X_15255_ _15255_/A _15277_/B vssd1 vssd1 vccd1 vccd1 _15263_/B sky130_fd_sc_hd__nor2_2
XFILLER_172_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12467_ _12465_/Y _12467_/B _12467_/C vssd1 vssd1 vccd1 vccd1 _12468_/A sky130_fd_sc_hd__and3b_1
X_14206_ _14206_/A _14330_/B vssd1 vssd1 vccd1 vccd1 _14206_/Y sky130_fd_sc_hd__nor2_1
XFILLER_125_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11418_ _17880_/Q vssd1 vssd1 vccd1 vccd1 _12316_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_193_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15186_ _15220_/A _15186_/B _15199_/C vssd1 vssd1 vccd1 vccd1 _15186_/X sky130_fd_sc_hd__or3_1
X_12398_ _12406_/B _12398_/B _12490_/A vssd1 vssd1 vccd1 vccd1 _12399_/A sky130_fd_sc_hd__and3b_1
XFILLER_67_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14137_ _18362_/Q _13562_/A _13568_/A _18356_/Q _14136_/X vssd1 vssd1 vccd1 vccd1
+ _14137_/X sky130_fd_sc_hd__a221o_1
XFILLER_119_1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11349_ _11357_/B vssd1 vssd1 vccd1 vccd1 _11495_/B sky130_fd_sc_hd__buf_2
XFILLER_67_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14068_ _18824_/Q _13581_/X _13582_/X _18818_/Q _14067_/X vssd1 vssd1 vccd1 vccd1
+ _14068_/X sky130_fd_sc_hd__a221o_1
X_18945_ _18950_/CLK _18945_/D vssd1 vssd1 vccd1 vccd1 _18945_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_98_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13019_ _18151_/Q _13019_/B vssd1 vssd1 vccd1 vccd1 _13039_/B sky130_fd_sc_hd__and2_1
XFILLER_80_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18876_ _18914_/CLK _18876_/D vssd1 vssd1 vccd1 vccd1 _18876_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_230_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17827_ _18157_/CLK _17827_/D vssd1 vssd1 vccd1 vccd1 _17827_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_54_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_214_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17758_ _17764_/A _19023_/Q vssd1 vssd1 vccd1 vccd1 _17759_/A sky130_fd_sc_hd__and2_1
XFILLER_81_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16709_ _16712_/B _16706_/X _16708_/Y _16704_/X vssd1 vssd1 vccd1 vccd1 _18745_/D
+ sky130_fd_sc_hd__o211a_1
X_17689_ _14597_/A _17687_/Y _17675_/X _17688_/Y _18984_/Q vssd1 vssd1 vccd1 vccd1
+ _17690_/B sky130_fd_sc_hd__a32o_1
XFILLER_165_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_222_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_200_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_222_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_200_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09112_ _18752_/Q _18751_/Q _18750_/Q vssd1 vssd1 vccd1 vccd1 _09114_/C sky130_fd_sc_hd__or3_4
Xclkbuf_leaf_152_wb_clk_i _18102_/CLK vssd1 vssd1 vccd1 vccd1 _18130_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_206_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09043_ _09046_/A vssd1 vssd1 vccd1 vccd1 _09043_/Y sky130_fd_sc_hd__inv_2
XFILLER_163_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_135_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_191_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_1238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09945_ _10307_/S vssd1 vssd1 vccd1 vccd1 _09945_/X sky130_fd_sc_hd__buf_6
XFILLER_213_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09876_ _09876_/A _09876_/B vssd1 vssd1 vccd1 vccd1 _09896_/B sky130_fd_sc_hd__xor2_2
XFILLER_112_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_213_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_12 _10722_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_23 _09243_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_34 _09924_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_45 _10403_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_56 _12285_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_67 _13734_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINSDIODE2_78 _13561_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_89 _13663_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_226_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_183_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10720_ _09153_/A _09143_/B _10841_/A vssd1 vssd1 vccd1 vccd1 _10720_/X sky130_fd_sc_hd__mux2_1
XFILLER_54_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10651_ _10779_/A vssd1 vssd1 vccd1 vccd1 _10805_/A sky130_fd_sc_hd__buf_2
XFILLER_224_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_220_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10582_ _10580_/X _10581_/X _10582_/S vssd1 vssd1 vccd1 vccd1 _10582_/X sky130_fd_sc_hd__mux2_1
X_13370_ _17768_/A _13370_/B _13370_/C vssd1 vssd1 vccd1 vccd1 _13371_/A sky130_fd_sc_hd__and3_1
XFILLER_221_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12321_ _17884_/Q _11431_/B _12316_/X vssd1 vssd1 vccd1 vccd1 _12327_/C sky130_fd_sc_hd__o21a_1
XFILLER_103_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15040_ _15184_/A _15085_/B vssd1 vssd1 vccd1 vccd1 _15049_/B sky130_fd_sc_hd__nor2_2
X_12252_ _11896_/X _12253_/A _12246_/Y _12250_/X _12251_/X vssd1 vssd1 vccd1 vccd1
+ _17862_/D sky130_fd_sc_hd__a41o_1
X_11203_ _11203_/A vssd1 vssd1 vccd1 vccd1 _17812_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_122_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12183_ _17849_/Q _12183_/B vssd1 vssd1 vccd1 vccd1 _12183_/X sky130_fd_sc_hd__and2_1
XFILLER_79_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_1305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11134_ _11595_/A vssd1 vssd1 vccd1 vccd1 _11582_/A sky130_fd_sc_hd__buf_2
XFILLER_1_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16991_ _18846_/Q _18810_/Q _17005_/S vssd1 vssd1 vccd1 vccd1 _16991_/X sky130_fd_sc_hd__mux2_1
XFILLER_122_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_231_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15942_ _15942_/A _15942_/B vssd1 vssd1 vccd1 vccd1 _15942_/Y sky130_fd_sc_hd__nand2_1
X_18730_ _18765_/CLK _18730_/D vssd1 vssd1 vccd1 vccd1 _18730_/Q sky130_fd_sc_hd__dfxtp_1
X_11065_ _17788_/Q vssd1 vssd1 vccd1 vccd1 _11942_/A sky130_fd_sc_hd__buf_4
XTAP_5230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_231_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10016_ _09153_/D _09148_/D _10019_/S vssd1 vssd1 vccd1 vccd1 _10016_/X sky130_fd_sc_hd__mux2_1
XTAP_5274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18661_ _18696_/CLK _18661_/D vssd1 vssd1 vccd1 vccd1 _18661_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_37_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15873_ _15873_/A _15876_/B vssd1 vssd1 vccd1 vccd1 _15873_/Y sky130_fd_sc_hd__nand2_1
XTAP_4540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14824_ _14827_/B _14821_/X _14823_/Y _14819_/X vssd1 vssd1 vccd1 vccd1 _18295_/D
+ sky130_fd_sc_hd__o211a_1
X_17612_ _17640_/A vssd1 vssd1 vccd1 vccd1 _17638_/A sky130_fd_sc_hd__clkbuf_1
X_18592_ _18593_/CLK _18592_/D vssd1 vssd1 vccd1 vccd1 _18592_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_229_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_205_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17543_ _18986_/Q _18950_/Q _17543_/S vssd1 vssd1 vccd1 vccd1 _17543_/X sky130_fd_sc_hd__mux2_1
XTAP_3883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14755_ _15197_/A _14790_/B vssd1 vssd1 vccd1 vccd1 _14767_/B sky130_fd_sc_hd__nor2_2
XTAP_3894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11967_ _11967_/A _13434_/B vssd1 vssd1 vccd1 vccd1 _12044_/A sky130_fd_sc_hd__nor2_1
XFILLER_17_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13706_ _13706_/A vssd1 vssd1 vccd1 vccd1 _13706_/X sky130_fd_sc_hd__buf_6
XFILLER_204_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17474_ _18930_/Q _17477_/B _17473_/X _17461_/X vssd1 vssd1 vccd1 vccd1 _18930_/D
+ sky130_fd_sc_hd__o211a_1
X_10918_ _10914_/X _10917_/X _10918_/S vssd1 vssd1 vccd1 vccd1 _10918_/X sky130_fd_sc_hd__mux2_1
XFILLER_229_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_220_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14686_ _16959_/A vssd1 vssd1 vccd1 vccd1 _15277_/A sky130_fd_sc_hd__buf_6
XFILLER_205_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11898_ _11209_/A _11896_/X _11011_/C _11897_/X vssd1 vssd1 vccd1 vccd1 _17838_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_60_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16425_ _18712_/Q _18676_/Q _16449_/S vssd1 vssd1 vccd1 vccd1 _16425_/X sky130_fd_sc_hd__mux2_1
XFILLER_20_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19213_ _19213_/A _08965_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[13] sky130_fd_sc_hd__ebufn_8
XFILLER_204_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13637_ _13710_/A _13637_/B vssd1 vssd1 vccd1 vccd1 _13637_/Y sky130_fd_sc_hd__nor2_2
XFILLER_220_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10849_ _10733_/X _10774_/X _10822_/X _10833_/X _10848_/X vssd1 vssd1 vccd1 vccd1
+ _10849_/X sky130_fd_sc_hd__a2111o_1
X_19144_ _19144_/A _09050_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[14] sky130_fd_sc_hd__ebufn_8
X_16356_ _16794_/A _16356_/B vssd1 vssd1 vccd1 vccd1 _16364_/B sky130_fd_sc_hd__nor2_1
X_13568_ _13568_/A vssd1 vssd1 vccd1 vccd1 _13568_/X sky130_fd_sc_hd__buf_4
XFILLER_160_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15307_ _18146_/Q _15772_/B vssd1 vssd1 vccd1 vccd1 _15440_/A sky130_fd_sc_hd__nand2_4
XFILLER_146_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_121_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12519_ _11767_/A _17427_/S _12514_/A _11769_/X vssd1 vssd1 vccd1 vccd1 _12520_/B
+ sky130_fd_sc_hd__o2bb2a_1
X_16287_ _16287_/A _16358_/C vssd1 vssd1 vccd1 vccd1 _16294_/B sky130_fd_sc_hd__nor2_2
XFILLER_200_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_185_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13499_ _13592_/A vssd1 vssd1 vccd1 vccd1 _13500_/A sky130_fd_sc_hd__buf_6
XFILLER_67_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18026_ _18030_/CLK _18026_/D vssd1 vssd1 vccd1 vccd1 _18026_/Q sky130_fd_sc_hd__dfxtp_1
X_15238_ _18434_/Q _18398_/Q _15246_/S vssd1 vssd1 vccd1 vccd1 _15238_/X sky130_fd_sc_hd__mux2_1
Xclkbuf_3_2_0_wb_clk_i clkbuf_3_3_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_4_5_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_2
X_15169_ _15182_/A _15169_/B vssd1 vssd1 vccd1 vccd1 _15169_/Y sky130_fd_sc_hd__nand2_1
XFILLER_160_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09730_ _17783_/Q vssd1 vssd1 vccd1 vccd1 _09742_/A sky130_fd_sc_hd__clkbuf_2
X_18928_ _18939_/CLK _18928_/D vssd1 vssd1 vccd1 vccd1 _18928_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_39_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_227_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09661_ _10204_/A _10623_/A vssd1 vssd1 vccd1 vccd1 _09661_/X sky130_fd_sc_hd__and2_1
XFILLER_228_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18859_ _18860_/CLK _18859_/D vssd1 vssd1 vccd1 vccd1 _18859_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_94_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_228_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09592_ _09598_/S _09592_/B vssd1 vssd1 vccd1 vccd1 _09593_/C sky130_fd_sc_hd__xor2_1
XFILLER_215_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_224_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_223_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_160 _18357_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINSDIODE2_171 _18856_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_182 _08972_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_193 _09143_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_206_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_1302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_1207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09026_ _09028_/A vssd1 vssd1 vccd1 vccd1 _09026_/Y sky130_fd_sc_hd__inv_2
XFILLER_108_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_176_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19085__56 vssd1 vssd1 vccd1 vccd1 _19085__56/HI _19193_/A sky130_fd_sc_hd__conb_1
X_09928_ _09392_/C _09397_/B _09402_/D _09397_/D _09909_/X _12121_/A vssd1 vssd1 vccd1
+ vccd1 _09928_/X sky130_fd_sc_hd__mux4_1
XFILLER_120_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_219_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_213_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09859_ _09879_/A _09879_/B vssd1 vssd1 vccd1 vccd1 _09860_/C sky130_fd_sc_hd__nor2_1
XFILLER_59_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_213_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12870_ _17953_/Q _12868_/B _12871_/B _12862_/X vssd1 vssd1 vccd1 vccd1 _17953_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_3135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11821_ _12257_/A vssd1 vssd1 vccd1 vccd1 _17556_/A sky130_fd_sc_hd__buf_8
XTAP_2434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_214_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14540_ _18232_/Q _14545_/B _14539_/Y _14533_/X vssd1 vssd1 vccd1 vccd1 _18232_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_1733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11752_ _11729_/X _11730_/Y _11750_/Y _11856_/C vssd1 vssd1 vccd1 vccd1 _11752_/X
+ sky130_fd_sc_hd__a211o_1
XTAP_1744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10703_ _09203_/A _09198_/C _09193_/D _09203_/D _10856_/S _10680_/A vssd1 vssd1 vccd1
+ vccd1 _10703_/X sky130_fd_sc_hd__mux4_2
XTAP_1777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14471_ _14504_/B _14471_/B _14471_/C vssd1 vssd1 vccd1 vccd1 _14472_/A sky130_fd_sc_hd__and3_1
XTAP_1788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11683_ _11683_/A _11683_/B _11683_/C vssd1 vssd1 vccd1 vccd1 _11683_/X sky130_fd_sc_hd__and3_1
XFILLER_14_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_197_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16210_ _16217_/B _16206_/X _16208_/X _16209_/X vssd1 vssd1 vccd1 vccd1 _18624_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_224_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13422_ _13442_/B vssd1 vssd1 vccd1 vccd1 _13422_/Y sky130_fd_sc_hd__inv_2
XFILLER_201_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10634_ _10838_/A vssd1 vssd1 vccd1 vccd1 _10864_/A sky130_fd_sc_hd__buf_2
X_17190_ _18860_/Q _17189_/B _17189_/Y _17181_/X vssd1 vssd1 vccd1 vccd1 _18860_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_220_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16141_ _18646_/Q _18610_/Q _16145_/S vssd1 vssd1 vccd1 vccd1 _16141_/X sky130_fd_sc_hd__mux2_1
XFILLER_195_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13353_ _13353_/A _13389_/B vssd1 vssd1 vccd1 vccd1 _13353_/Y sky130_fd_sc_hd__nand2_1
X_10565_ _10903_/S _10558_/Y _10564_/Y _10533_/B _10547_/A vssd1 vssd1 vccd1 vccd1
+ _10897_/A sky130_fd_sc_hd__a2111oi_1
XFILLER_182_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12304_ _12304_/A _12304_/B _12327_/B vssd1 vssd1 vccd1 vccd1 _12304_/Y sky130_fd_sc_hd__nor3_1
X_16072_ _16823_/A vssd1 vssd1 vccd1 vccd1 _16678_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_143_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13284_ _18033_/Q _18032_/Q _18035_/Q _18034_/Q vssd1 vssd1 vccd1 vccd1 _13286_/C
+ sky130_fd_sc_hd__or4_1
X_10496_ _10496_/A _10496_/B vssd1 vssd1 vccd1 vccd1 _10496_/Y sky130_fd_sc_hd__nand2_1
XFILLER_136_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15023_ _15025_/B _15021_/X _15022_/Y _15004_/X vssd1 vssd1 vccd1 vccd1 _18343_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_142_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12235_ _12235_/A _12239_/C vssd1 vssd1 vccd1 vccd1 _12235_/Y sky130_fd_sc_hd__nor2_1
XFILLER_216_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_122_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12166_ _17844_/Q _12172_/B _12165_/Y vssd1 vssd1 vccd1 vccd1 _12166_/X sky130_fd_sc_hd__a21o_1
XFILLER_2_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11117_ _11452_/A vssd1 vssd1 vccd1 vccd1 _11788_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_190_1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_231_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16974_ _17412_/A vssd1 vssd1 vccd1 vccd1 _16975_/A sky130_fd_sc_hd__buf_2
X_12097_ _13526_/C _12097_/B vssd1 vssd1 vccd1 vccd1 _12104_/B sky130_fd_sc_hd__xnor2_1
XFILLER_1_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18713_ _18719_/CLK _18713_/D vssd1 vssd1 vccd1 vccd1 _18713_/Q sky130_fd_sc_hd__dfxtp_4
X_15925_ _15925_/A vssd1 vssd1 vccd1 vccd1 _15925_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_209_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11048_ _13375_/A _17997_/Q _17996_/Q _13394_/D vssd1 vssd1 vccd1 vccd1 _13383_/A
+ sky130_fd_sc_hd__and4bb_4
XTAP_5071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18644_ _18668_/CLK _18644_/D vssd1 vssd1 vccd1 vccd1 _18644_/Q sky130_fd_sc_hd__dfxtp_2
X_15856_ _18579_/Q _18543_/Q _15859_/S vssd1 vssd1 vccd1 vccd1 _15856_/X sky130_fd_sc_hd__mux2_1
XFILLER_37_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14807_ _14856_/A _15243_/B _14818_/C vssd1 vssd1 vccd1 vccd1 _14807_/X sky130_fd_sc_hd__or3_1
XFILLER_64_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_206_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15787_ _18561_/Q _18525_/Q _15790_/S vssd1 vssd1 vccd1 vccd1 _15787_/X sky130_fd_sc_hd__mux2_1
X_18575_ _18577_/CLK _18575_/D vssd1 vssd1 vccd1 vccd1 _18575_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_75_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12999_ _13000_/B _12990_/A _13000_/A vssd1 vssd1 vccd1 vccd1 _13001_/A sky130_fd_sc_hd__a21oi_1
XFILLER_51_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_1351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14738_ _14778_/A vssd1 vssd1 vccd1 vccd1 _14738_/X sky130_fd_sc_hd__clkbuf_2
X_17526_ _17526_/A _17536_/B vssd1 vssd1 vccd1 vccd1 _17534_/B sky130_fd_sc_hd__nor2_1
XFILLER_32_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_220_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17457_ _17456_/B _17455_/X _17456_/Y _17441_/X vssd1 vssd1 vccd1 vccd1 _18926_/D
+ sky130_fd_sc_hd__o211a_1
X_14669_ _18259_/Q _14670_/B _14667_/Y _14668_/X vssd1 vssd1 vccd1 vccd1 _18259_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_221_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_220_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16408_ _16407_/B _16405_/X _16407_/Y _16398_/X vssd1 vssd1 vccd1 vccd1 _18671_/D
+ sky130_fd_sc_hd__o211a_1
X_17388_ _17437_/A _17528_/B _17399_/C vssd1 vssd1 vccd1 vccd1 _17388_/X sky130_fd_sc_hd__or3_1
XFILLER_146_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_220_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_203_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16339_ _16342_/B _16336_/X _16338_/Y _16334_/X vssd1 vssd1 vccd1 vccd1 _18655_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_9_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_203_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_1240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_1330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18009_ _18213_/CLK _18009_/D vssd1 vssd1 vccd1 vccd1 _18009_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_86_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_1333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_142_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09713_ _18257_/Q _18256_/Q _18255_/Q vssd1 vssd1 vccd1 vccd1 _09713_/X sky130_fd_sc_hd__or3_4
XFILLER_210_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_216_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09644_ _13353_/A vssd1 vssd1 vccd1 vccd1 _09647_/A sky130_fd_sc_hd__inv_2
XFILLER_216_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_222_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_215_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09575_ _09575_/A _09575_/B vssd1 vssd1 vccd1 vccd1 _09585_/A sky130_fd_sc_hd__nor2_1
XFILLER_93_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_224_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_223_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_196_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_221_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_221_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_192_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10350_ _10350_/A _10391_/B vssd1 vssd1 vccd1 vccd1 _10350_/X sky130_fd_sc_hd__or2_1
XFILLER_109_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09009_ _09010_/A vssd1 vssd1 vccd1 vccd1 _09009_/Y sky130_fd_sc_hd__inv_2
XFILLER_178_1288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10281_ _10281_/A _10281_/B vssd1 vssd1 vccd1 vccd1 _10281_/Y sky130_fd_sc_hd__nor2_1
XFILLER_2_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12020_ _12020_/A _12020_/B vssd1 vssd1 vccd1 vccd1 _12022_/C sky130_fd_sc_hd__and2_4
XFILLER_183_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13971_ _18283_/Q _13666_/X _13624_/A _18277_/Q vssd1 vssd1 vccd1 vccd1 _13971_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_65_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15710_ _16005_/A _15745_/B vssd1 vssd1 vccd1 vccd1 _15719_/B sky130_fd_sc_hd__nor2_1
XFILLER_19_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12922_ _12956_/A vssd1 vssd1 vccd1 vccd1 _12983_/A sky130_fd_sc_hd__buf_2
X_16690_ _18777_/Q _18741_/Q _16694_/S vssd1 vssd1 vccd1 vccd1 _16690_/X sky130_fd_sc_hd__mux2_1
XFILLER_18_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15641_ _15651_/B _15637_/X _15638_/X _15640_/X vssd1 vssd1 vccd1 vccd1 _18489_/D
+ sky130_fd_sc_hd__o211a_1
X_12853_ _12853_/A vssd1 vssd1 vccd1 vccd1 _17948_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18360_ _18367_/CLK _18360_/D vssd1 vssd1 vccd1 vccd1 _18360_/Q sky130_fd_sc_hd__dfxtp_2
X_11804_ _11976_/A _11976_/B vssd1 vssd1 vccd1 vccd1 _11964_/A sky130_fd_sc_hd__nand2_2
XFILLER_73_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15572_ _16019_/A _15597_/B vssd1 vssd1 vccd1 vccd1 _15583_/B sky130_fd_sc_hd__nor2_2
XTAP_1530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12784_ _13080_/A _12784_/B _13066_/C vssd1 vssd1 vccd1 vccd1 _12784_/X sky130_fd_sc_hd__or3_1
XTAP_2275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17311_ _17334_/A _17314_/B vssd1 vssd1 vccd1 vccd1 _17311_/Y sky130_fd_sc_hd__nand2_1
XFILLER_230_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_202_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14523_ _14702_/A vssd1 vssd1 vccd1 vccd1 _17415_/B sky130_fd_sc_hd__clkbuf_8
XPHY_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18291_ _18312_/CLK _18291_/D vssd1 vssd1 vccd1 vccd1 _18291_/Q sky130_fd_sc_hd__dfxtp_1
X_11735_ _11735_/A _11735_/B vssd1 vssd1 vccd1 vccd1 _11740_/B sky130_fd_sc_hd__or2_1
XPHY_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17242_ _17240_/B _17239_/X _17240_/Y _17241_/X vssd1 vssd1 vccd1 vccd1 _18872_/D
+ sky130_fd_sc_hd__o211a_1
X_14454_ _18204_/Q _14453_/X _14428_/X _09506_/B vssd1 vssd1 vccd1 vccd1 _14455_/B
+ sky130_fd_sc_hd__o2bb2a_1
X_11666_ _11639_/A _11651_/A _11668_/A vssd1 vssd1 vccd1 vccd1 _11666_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_128_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13405_ _17768_/A _13405_/B _13405_/C vssd1 vssd1 vccd1 vccd1 _13406_/A sky130_fd_sc_hd__and3_1
XFILLER_179_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10617_ _10675_/A vssd1 vssd1 vccd1 vccd1 _13007_/A sky130_fd_sc_hd__clkbuf_4
X_17173_ _17193_/A _17460_/B _17173_/C vssd1 vssd1 vccd1 vccd1 _17173_/X sky130_fd_sc_hd__or3_1
X_14385_ _14399_/A vssd1 vssd1 vccd1 vccd1 _14386_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_167_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11597_ _11764_/A _11635_/A _11597_/C vssd1 vssd1 vccd1 vccd1 _11598_/B sky130_fd_sc_hd__or3_1
X_16124_ _16123_/B _16122_/X _16123_/Y _16120_/X vssd1 vssd1 vccd1 vccd1 _18605_/D
+ sky130_fd_sc_hd__o211a_1
X_13336_ _13344_/A vssd1 vssd1 vccd1 vccd1 _13336_/X sky130_fd_sc_hd__clkbuf_2
X_10548_ _09198_/A _09193_/A _09203_/B _10293_/A _10521_/A _10550_/S vssd1 vssd1 vccd1
+ vccd1 _10549_/B sky130_fd_sc_hd__mux4_1
XFILLER_6_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16055_ _16055_/A _16208_/C vssd1 vssd1 vccd1 vccd1 _16064_/B sky130_fd_sc_hd__nor2_2
XFILLER_143_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13267_ _13267_/A vssd1 vssd1 vccd1 vccd1 _18086_/D sky130_fd_sc_hd__clkbuf_1
X_10479_ _09265_/C _09265_/A _09270_/A _10813_/A _10412_/A _10411_/A vssd1 vssd1 vccd1
+ vccd1 _10479_/X sky130_fd_sc_hd__mux4_1
XFILLER_142_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15006_ _15643_/A vssd1 vssd1 vccd1 vccd1 _15247_/A sky130_fd_sc_hd__clkbuf_2
X_12218_ _17747_/A vssd1 vssd1 vccd1 vccd1 _13037_/A sky130_fd_sc_hd__buf_2
XFILLER_68_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13198_ _13198_/A vssd1 vssd1 vccd1 vccd1 _18055_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_111_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12149_ _17840_/Q _12171_/B _12180_/B _11863_/X vssd1 vssd1 vccd1 vccd1 _17840_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_229_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16957_ _16957_/A _16957_/B vssd1 vssd1 vccd1 vccd1 _16957_/Y sky130_fd_sc_hd__nand2_1
XFILLER_81_1293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15908_ _16041_/B vssd1 vssd1 vccd1 vccd1 _15964_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_38_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16888_ _18825_/Q _18789_/Q _16900_/S vssd1 vssd1 vccd1 vccd1 _16888_/X sky130_fd_sc_hd__mux2_1
XFILLER_37_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18627_ _18650_/CLK _18627_/D vssd1 vssd1 vccd1 vccd1 _18627_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_64_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_225_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15839_ _15876_/A _15839_/B vssd1 vssd1 vccd1 vccd1 _15839_/Y sky130_fd_sc_hd__nand2_1
XFILLER_25_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09360_ _09360_/A _09360_/B _09360_/C _09360_/D vssd1 vssd1 vccd1 vccd1 _09371_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_80_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18558_ _18572_/CLK _18558_/D vssd1 vssd1 vccd1 vccd1 _18558_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_178_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_5_23_0_wb_clk_i clkbuf_5_23_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_5_23_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_162_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17509_ _17509_/A _17512_/B vssd1 vssd1 vccd1 vccd1 _17509_/Y sky130_fd_sc_hd__nand2_1
XFILLER_177_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09291_ _18491_/Q _18490_/Q _18489_/Q vssd1 vssd1 vccd1 vccd1 _09294_/B sky130_fd_sc_hd__or3_2
XFILLER_166_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18489_ _18497_/CLK _18489_/D vssd1 vssd1 vccd1 vccd1 _18489_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_178_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_220_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_177_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_59_wb_clk_i _18759_/CLK vssd1 vssd1 vccd1 vccd1 _18738_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_20_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_115_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19055__26 vssd1 vssd1 vccd1 vccd1 _19055__26/HI _19149_/A sky130_fd_sc_hd__conb_1
XFILLER_60_1322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_229_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_229_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_210_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_228_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_216_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_210_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09627_ _10204_/A _10629_/A vssd1 vssd1 vccd1 vccd1 _09627_/X sky130_fd_sc_hd__and2_1
XFILLER_216_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_1271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_231_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_1240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09558_ _12066_/A _12065_/A vssd1 vssd1 vccd1 vccd1 _10044_/A sky130_fd_sc_hd__and2_2
XFILLER_102_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09489_ _14507_/B vssd1 vssd1 vccd1 vccd1 _13416_/A sky130_fd_sc_hd__buf_6
XFILLER_145_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_200_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11520_ _11622_/A _11516_/X _11519_/X vssd1 vssd1 vccd1 vccd1 _11520_/X sky130_fd_sc_hd__a21o_1
XFILLER_184_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11451_ _11488_/A _11451_/B vssd1 vssd1 vccd1 vccd1 _11451_/Y sky130_fd_sc_hd__nor2_1
XFILLER_11_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_221_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10402_ _09895_/X _10400_/X _10401_/X _10278_/X vssd1 vssd1 vccd1 vccd1 _10403_/B
+ sky130_fd_sc_hd__a22oi_4
XFILLER_183_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14170_ _18611_/Q _14124_/X _13538_/A _18593_/Q vssd1 vssd1 vccd1 vccd1 _14170_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_164_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11382_ _11525_/B vssd1 vssd1 vccd1 vccd1 _11619_/A sky130_fd_sc_hd__buf_2
XFILLER_3_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13121_ _13129_/A _18021_/Q vssd1 vssd1 vccd1 vccd1 _13122_/A sky130_fd_sc_hd__and2_1
X_10333_ _10331_/X _10332_/X _10333_/S vssd1 vssd1 vccd1 vccd1 _10333_/X sky130_fd_sc_hd__mux2_1
XFILLER_125_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13052_ _18002_/Q _18004_/Q _13058_/B vssd1 vssd1 vccd1 vccd1 _13052_/X sky130_fd_sc_hd__and3_1
XFILLER_191_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10264_ _10264_/A _10264_/B vssd1 vssd1 vccd1 vccd1 _10513_/A sky130_fd_sc_hd__xnor2_4
XFILLER_3_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12003_ _12007_/A _12020_/B _12021_/B vssd1 vssd1 vccd1 vccd1 _12043_/A sky130_fd_sc_hd__o21ai_1
XFILLER_152_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17860_ _19035_/CLK _17860_/D vssd1 vssd1 vccd1 vccd1 _17860_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_78_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10195_ _18099_/Q _12946_/A vssd1 vssd1 vccd1 vccd1 _10195_/X sky130_fd_sc_hd__and2_1
XFILLER_152_1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16811_ _16866_/A _17415_/B _16866_/C vssd1 vssd1 vccd1 vccd1 _16811_/X sky130_fd_sc_hd__or3_1
XFILLER_120_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17791_ _17793_/CLK _17791_/D vssd1 vssd1 vccd1 vccd1 _17791_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_120_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13954_ _18517_/Q _13730_/X _13732_/X _18508_/Q _13953_/X vssd1 vssd1 vccd1 vccd1
+ _13954_/X sky130_fd_sc_hd__a221o_2
X_16742_ _18791_/Q _18755_/Q _16742_/S vssd1 vssd1 vccd1 vccd1 _16742_/X sky130_fd_sc_hd__mux2_1
XFILLER_4_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12905_ _17963_/Q _17964_/Q _12899_/B _17965_/Q vssd1 vssd1 vccd1 vccd1 _12906_/C
+ sky130_fd_sc_hd__a31o_1
X_16673_ _16673_/A vssd1 vssd1 vccd1 vccd1 _17278_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_62_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13885_ _18973_/Q _13848_/A _13877_/A _18967_/Q _13884_/X vssd1 vssd1 vccd1 vccd1
+ _13885_/X sky130_fd_sc_hd__a221o_1
XFILLER_185_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18412_ _18432_/CLK _18412_/D vssd1 vssd1 vccd1 vccd1 _18412_/Q sky130_fd_sc_hd__dfxtp_1
X_15624_ _18522_/Q _18486_/Q _15642_/S vssd1 vssd1 vccd1 vccd1 _15624_/X sky130_fd_sc_hd__mux2_1
XFILLER_34_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12836_ _12814_/X _12823_/X _12835_/X _12361_/A vssd1 vssd1 vccd1 vccd1 _12847_/A
+ sky130_fd_sc_hd__o31a_1
XTAP_2050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_222_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_185_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_1310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15555_ _15616_/A vssd1 vssd1 vccd1 vccd1 _15555_/X sky130_fd_sc_hd__clkbuf_2
X_18343_ _18343_/CLK _18343_/D vssd1 vssd1 vccd1 vccd1 _18343_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_2094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_159_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12767_ _12775_/A vssd1 vssd1 vccd1 vccd1 _13269_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_203_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_202_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14506_ _14373_/A _14422_/A _14372_/B vssd1 vssd1 vccd1 vccd1 _14508_/A sky130_fd_sc_hd__a21oi_1
XFILLER_202_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18274_ _18278_/CLK _18274_/D vssd1 vssd1 vccd1 vccd1 _18274_/Q sky130_fd_sc_hd__dfxtp_1
X_11718_ _17912_/Q vssd1 vssd1 vccd1 vccd1 _11720_/A sky130_fd_sc_hd__inv_2
X_15486_ _18488_/Q _18452_/Q _15494_/S vssd1 vssd1 vccd1 vccd1 _15486_/X sky130_fd_sc_hd__mux2_1
XFILLER_175_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_1349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12698_ _12698_/A _12707_/B vssd1 vssd1 vccd1 vccd1 _12698_/Y sky130_fd_sc_hd__nor2_1
XFILLER_159_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14437_ _14434_/Y _14435_/X _14436_/X vssd1 vssd1 vccd1 vccd1 _18199_/D sky130_fd_sc_hd__o21a_1
X_17225_ _17230_/B _17221_/X _17224_/Y _17219_/X vssd1 vssd1 vccd1 vccd1 _18868_/D
+ sky130_fd_sc_hd__o211a_1
X_11649_ _12251_/A _11648_/X _11339_/B _11639_/A vssd1 vssd1 vccd1 vccd1 _11649_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_156_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_174_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17156_ _17156_/A _17156_/B vssd1 vssd1 vccd1 vccd1 _17156_/Y sky130_fd_sc_hd__nand2_1
X_14368_ _18185_/Q _14366_/Y _14367_/X _14340_/X vssd1 vssd1 vccd1 vccd1 _18185_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_155_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_200_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16107_ _16109_/B _16105_/X _16106_/Y _16097_/X vssd1 vssd1 vccd1 vccd1 _18601_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_115_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13319_ _13322_/B _13317_/Y _13318_/X vssd1 vssd1 vccd1 vccd1 _13319_/X sky130_fd_sc_hd__a21o_1
X_17087_ _18871_/Q _18835_/Q _17094_/S vssd1 vssd1 vccd1 vccd1 _17087_/X sky130_fd_sc_hd__mux2_1
XFILLER_115_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14299_ _14299_/A vssd1 vssd1 vccd1 vccd1 _14299_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_171_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16038_ _18623_/Q _18587_/Q _16050_/S vssd1 vssd1 vccd1 vccd1 _16038_/X sky130_fd_sc_hd__mux2_1
XFILLER_157_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_1366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_177_wb_clk_i clkbuf_5_11_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18224_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_69_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_106_wb_clk_i clkbuf_5_29_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18542_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_170_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17989_ _18044_/CLK _17989_/D vssd1 vssd1 vccd1 vccd1 _17989_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_85_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_111_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_1366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09412_ _18320_/Q _18319_/Q _18318_/Q vssd1 vssd1 vccd1 vccd1 _09413_/D sky130_fd_sc_hd__or3_2
XFILLER_53_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_1298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09343_ _18422_/Q _18421_/Q _18420_/Q vssd1 vssd1 vccd1 vccd1 _09344_/D sky130_fd_sc_hd__or3_4
XFILLER_12_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_1348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_178_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09274_ _18875_/Q _18874_/Q _18873_/Q vssd1 vssd1 vccd1 vccd1 _09277_/B sky130_fd_sc_hd__or3_2
XFILLER_20_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_148_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_1271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_147_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_134_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_138_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08989_ _08991_/A vssd1 vssd1 vccd1 vccd1 _08989_/Y sky130_fd_sc_hd__inv_2
XTAP_5659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_229_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_91_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_216_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10951_ _09402_/A _09392_/B _09397_/C _10877_/A _10003_/S _09987_/X vssd1 vssd1 vccd1
+ vccd1 _10952_/B sky130_fd_sc_hd__mux4_1
XFILLER_44_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_216_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13670_ _13670_/A vssd1 vssd1 vccd1 vccd1 _13670_/X sky130_fd_sc_hd__buf_6
XFILLER_44_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10882_ _09365_/A _09370_/B _10882_/S vssd1 vssd1 vccd1 vccd1 _10882_/X sky130_fd_sc_hd__mux2_1
XFILLER_16_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12621_ _12708_/A vssd1 vssd1 vccd1 vccd1 _12621_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_71_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15340_ _15404_/A vssd1 vssd1 vccd1 vccd1 _15340_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_12_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12552_ _12588_/B _12809_/A vssd1 vssd1 vccd1 vccd1 _12554_/A sky130_fd_sc_hd__nor2_1
XFILLER_200_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11503_ _11503_/A _11719_/B vssd1 vssd1 vccd1 vccd1 _11742_/A sky130_fd_sc_hd__nor2_2
X_15271_ _18442_/Q _18406_/Q _15285_/S vssd1 vssd1 vccd1 vccd1 _15271_/X sky130_fd_sc_hd__mux2_1
X_12483_ _12480_/Y _12484_/B _12482_/X vssd1 vssd1 vccd1 vccd1 _17908_/D sky130_fd_sc_hd__a21boi_1
XFILLER_12_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17010_ _17035_/A _17010_/B vssd1 vssd1 vccd1 vccd1 _17010_/Y sky130_fd_sc_hd__nand2_1
X_14222_ _14222_/A _14305_/A vssd1 vssd1 vccd1 vccd1 _14222_/Y sky130_fd_sc_hd__nor2_1
X_11434_ _11415_/Y _12329_/B _11433_/X _11428_/Y vssd1 vssd1 vccd1 vccd1 _11434_/X
+ sky130_fd_sc_hd__o31a_1
XFILLER_184_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14153_ _18740_/Q _13508_/A _13515_/A _18746_/Q vssd1 vssd1 vccd1 vccd1 _14153_/X
+ sky130_fd_sc_hd__a22o_1
X_11365_ _11547_/B _11365_/B _11790_/B _11468_/B vssd1 vssd1 vccd1 vccd1 _11843_/B
+ sky130_fd_sc_hd__or4_1
XFILLER_193_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_4_wb_clk_i _17929_/CLK vssd1 vssd1 vccd1 vccd1 _18991_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_98_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13104_ _13104_/A vssd1 vssd1 vccd1 vccd1 _18012_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_113_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10316_ _09270_/B _09260_/D _10316_/S vssd1 vssd1 vccd1 vccd1 _10316_/X sky130_fd_sc_hd__mux2_1
X_14084_ _18461_/Q _13493_/A _13861_/X _18476_/Q vssd1 vssd1 vccd1 vccd1 _14084_/X
+ sky130_fd_sc_hd__a22o_1
X_18961_ _18972_/CLK _18961_/D vssd1 vssd1 vccd1 vccd1 _18961_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_112_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11296_ _11334_/B _11312_/B vssd1 vssd1 vccd1 vccd1 _11296_/Y sky130_fd_sc_hd__nand2_1
XFILLER_98_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13035_ _17990_/Q _13015_/X _13034_/X vssd1 vssd1 vccd1 vccd1 _17990_/D sky130_fd_sc_hd__a21o_1
X_17912_ _18960_/CLK _17912_/D vssd1 vssd1 vccd1 vccd1 _17912_/Q sky130_fd_sc_hd__dfxtp_2
X_10247_ _18120_/Q vssd1 vssd1 vccd1 vccd1 _10253_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_18892_ _18893_/CLK _18892_/D vssd1 vssd1 vccd1 vccd1 _18892_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_224_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17843_ _19019_/CLK _17843_/D vssd1 vssd1 vccd1 vccd1 _17843_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10178_ _10178_/A _10178_/B vssd1 vssd1 vccd1 vccd1 _10179_/B sky130_fd_sc_hd__xnor2_2
XFILLER_113_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17774_ _11549_/X _12266_/X _12178_/X vssd1 vssd1 vccd1 vccd1 _19032_/D sky130_fd_sc_hd__o21a_1
XFILLER_66_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14986_ _18372_/Q _18336_/Q _14994_/S vssd1 vssd1 vccd1 vccd1 _14986_/X sky130_fd_sc_hd__mux2_1
XFILLER_130_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_219_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16725_ _16723_/B _16722_/X _16723_/Y _16724_/X vssd1 vssd1 vccd1 vccd1 _18749_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_19_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13937_ _18310_/Q _13749_/X _13933_/X _13936_/X vssd1 vssd1 vccd1 vccd1 _13937_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_208_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_208_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13868_ _18478_/Q _13617_/X _13619_/X _18454_/Q vssd1 vssd1 vccd1 vccd1 _13868_/X
+ sky130_fd_sc_hd__a22o_1
X_16656_ _16658_/B _16654_/X _16655_/Y _16639_/X vssd1 vssd1 vccd1 vccd1 _18733_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_37_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12819_ _17955_/Q vssd1 vssd1 vccd1 vccd1 _12824_/A sky130_fd_sc_hd__clkbuf_2
X_15607_ _15463_/B _15607_/B _15607_/C vssd1 vssd1 vccd1 vccd1 _17410_/A sky130_fd_sc_hd__nand3b_4
XFILLER_90_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_222_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13799_ _18360_/Q _13716_/X _13579_/A _18354_/Q _13798_/X vssd1 vssd1 vccd1 vccd1
+ _13799_/X sky130_fd_sc_hd__a221o_1
X_16587_ _17228_/A vssd1 vssd1 vccd1 vccd1 _16832_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_16_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18326_ _18350_/CLK _18326_/D vssd1 vssd1 vccd1 vccd1 _18326_/Q sky130_fd_sc_hd__dfxtp_4
X_15538_ _15982_/A _15548_/B vssd1 vssd1 vccd1 vccd1 _15546_/B sky130_fd_sc_hd__nor2_1
XFILLER_203_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15469_ _15492_/A _15909_/B _15515_/C vssd1 vssd1 vccd1 vccd1 _15469_/X sky130_fd_sc_hd__or3_1
X_18257_ _18266_/CLK _18257_/D vssd1 vssd1 vccd1 vccd1 _18257_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_191_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17208_ _17213_/B _17204_/X _17207_/X _17197_/X vssd1 vssd1 vccd1 vccd1 _18864_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_50_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_116_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18188_ _18230_/CLK _18188_/D vssd1 vssd1 vccd1 vccd1 _18188_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_156_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17139_ _17152_/A _17143_/B vssd1 vssd1 vccd1 vccd1 _17139_/Y sky130_fd_sc_hd__nand2_1
XFILLER_116_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09961_ _10598_/A vssd1 vssd1 vccd1 vccd1 _10388_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_171_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09892_ _09892_/A _09892_/B vssd1 vssd1 vccd1 vccd1 _09920_/B sky130_fd_sc_hd__xnor2_4
XFILLER_134_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_213_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_214_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_74_wb_clk_i clkbuf_5_21_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18683_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_222_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09326_ _18554_/Q _18553_/Q _18552_/Q vssd1 vssd1 vccd1 vccd1 _09327_/D sky130_fd_sc_hd__or3_4
XFILLER_16_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_1262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_181_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09257_ _18956_/Q _18955_/Q _18954_/Q vssd1 vssd1 vccd1 vccd1 _09260_/B sky130_fd_sc_hd__or3_4
XFILLER_21_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09188_ _09188_/A _09187_/Y vssd1 vssd1 vccd1 vccd1 _09188_/X sky130_fd_sc_hd__or2b_1
XFILLER_119_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_218_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_175_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_175_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11150_ _11150_/A vssd1 vssd1 vccd1 vccd1 _17802_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_122_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10101_ _09260_/A _09270_/C _09270_/D _09265_/D _09995_/A _09708_/A vssd1 vssd1 vccd1
+ vccd1 _10101_/X sky130_fd_sc_hd__mux4_1
XFILLER_108_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11081_ _11984_/C vssd1 vssd1 vccd1 vccd1 _11334_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_216_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_1364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10032_ _10012_/X _10031_/X _09728_/D vssd1 vssd1 vccd1 vccd1 _10032_/X sky130_fd_sc_hd__o21a_2
XTAP_5434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14840_ _14838_/B _14837_/X _14838_/Y _14839_/X vssd1 vssd1 vccd1 vccd1 _18299_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_75_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14771_ _17471_/A vssd1 vssd1 vccd1 vccd1 _15371_/B sky130_fd_sc_hd__buf_6
XFILLER_29_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_217_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11983_ _11983_/A _11983_/B vssd1 vssd1 vccd1 vccd1 _11985_/B sky130_fd_sc_hd__and2_1
XTAP_4799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16510_ _16510_/A _16510_/B vssd1 vssd1 vccd1 vccd1 _16510_/Y sky130_fd_sc_hd__nand2_1
X_13722_ _18234_/Q _13719_/X _13721_/X _18258_/Q vssd1 vssd1 vccd1 vccd1 _13722_/X
+ sky130_fd_sc_hd__a22o_1
Xclkbuf_4_4_0_wb_clk_i clkbuf_4_5_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_5_9_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_56_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10934_ _09304_/A _09294_/B _09299_/C _09304_/C _10495_/S _10522_/X vssd1 vssd1 vccd1
+ vccd1 _10934_/X sky130_fd_sc_hd__mux4_1
X_17490_ _17489_/B _17488_/X _17489_/Y _17478_/X vssd1 vssd1 vccd1 vccd1 _18935_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_17_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_216_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16441_ _16734_/A _16452_/B vssd1 vssd1 vccd1 vccd1 _16450_/B sky130_fd_sc_hd__nor2_2
XFILLER_182_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13653_ _13781_/A vssd1 vssd1 vccd1 vccd1 _13654_/A sky130_fd_sc_hd__buf_6
XFILLER_72_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10865_ _10600_/B _09676_/X _09677_/X _09678_/X _12092_/A _14206_/A vssd1 vssd1 vccd1
+ vccd1 _10865_/X sky130_fd_sc_hd__mux4_2
XFILLER_73_1321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_231_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12604_ _17925_/Q vssd1 vssd1 vccd1 vccd1 _12609_/B sky130_fd_sc_hd__clkbuf_2
X_16372_ _18663_/Q _16378_/B _16371_/X _16354_/X vssd1 vssd1 vccd1 vccd1 _18663_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_176_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19160_ _19160_/A _09024_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[30] sky130_fd_sc_hd__ebufn_8
X_13584_ _13760_/A vssd1 vssd1 vccd1 vccd1 _13585_/A sky130_fd_sc_hd__buf_6
XPHY_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10796_ _09214_/C _10687_/A _10795_/X _10770_/X vssd1 vssd1 vccd1 vccd1 _10796_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_223_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15323_ _15649_/A vssd1 vssd1 vccd1 vccd1 _15582_/A sky130_fd_sc_hd__clkbuf_2
XPHY_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18111_ _19028_/CLK _18111_/D vssd1 vssd1 vccd1 vccd1 _18111_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_158_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12535_ _12535_/A _12535_/B vssd1 vssd1 vccd1 vccd1 _12535_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_129_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_223_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_184_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15254_ _15253_/B _15251_/X _15253_/Y _15244_/X vssd1 vssd1 vccd1 vccd1 _18401_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_157_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18042_ _18094_/CLK _18042_/D vssd1 vssd1 vccd1 vccd1 _18042_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_201_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12466_ _12477_/C _12466_/B _12466_/C vssd1 vssd1 vccd1 vccd1 _12467_/B sky130_fd_sc_hd__nand3_1
XFILLER_173_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_144_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14205_ _14205_/A vssd1 vssd1 vccd1 vccd1 _14205_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_144_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11417_ _11423_/A vssd1 vssd1 vccd1 vccd1 _12329_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_15185_ _18420_/Q _18384_/Q _15198_/S vssd1 vssd1 vccd1 vccd1 _15185_/X sky130_fd_sc_hd__mux2_1
XFILLER_137_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12397_ _12397_/A _12397_/B _12397_/C vssd1 vssd1 vccd1 vccd1 _12398_/B sky130_fd_sc_hd__or3_1
XFILLER_193_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14136_ _18353_/Q _13492_/A _14030_/A _18368_/Q vssd1 vssd1 vccd1 vccd1 _14136_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_153_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11348_ _17795_/Q _11466_/B vssd1 vssd1 vccd1 vccd1 _11357_/B sky130_fd_sc_hd__and2_1
XFILLER_180_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_193_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14067_ _18830_/Q _13856_/A _13588_/X _18821_/Q vssd1 vssd1 vccd1 vccd1 _14067_/X
+ sky130_fd_sc_hd__a22o_1
X_18944_ _18953_/CLK _18944_/D vssd1 vssd1 vccd1 vccd1 _18944_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_113_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11279_ _17786_/Q _11333_/A _17787_/Q vssd1 vssd1 vccd1 vccd1 _13443_/A sky130_fd_sc_hd__o21a_1
XFILLER_79_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13018_ _17983_/Q _13015_/X _13017_/X vssd1 vssd1 vccd1 vccd1 _17983_/D sky130_fd_sc_hd__a21o_1
XFILLER_100_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_230_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18875_ _18875_/CLK _18875_/D vssd1 vssd1 vccd1 vccd1 _18875_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_227_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_228_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_230_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17826_ _18157_/CLK _17826_/D vssd1 vssd1 vccd1 vccd1 _17826_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_12_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17757_ _17757_/A vssd1 vssd1 vccd1 vccd1 _19021_/D sky130_fd_sc_hd__clkbuf_1
X_14969_ _14971_/B _14967_/X _14968_/Y _14961_/X vssd1 vssd1 vccd1 vccd1 _18331_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_47_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16708_ _16752_/A _16712_/B vssd1 vssd1 vccd1 vccd1 _16708_/Y sky130_fd_sc_hd__nand2_1
XFILLER_81_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17688_ _17687_/Y _17631_/A _14386_/A vssd1 vssd1 vccd1 vccd1 _17688_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_222_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16639_ _16659_/A vssd1 vssd1 vccd1 vccd1 _16639_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_165_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_223_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_222_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09111_ _18764_/Q _18763_/Q _18762_/Q vssd1 vssd1 vccd1 vccd1 _09114_/B sky130_fd_sc_hd__or3_4
X_18309_ _18312_/CLK _18309_/D vssd1 vssd1 vccd1 vccd1 _18309_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_202_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09042_ _09046_/A vssd1 vssd1 vccd1 vccd1 _09042_/Y sky130_fd_sc_hd__inv_2
XFILLER_108_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_191_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_209_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_192_wb_clk_i clkbuf_5_12_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18992_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_85_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_121_wb_clk_i clkbuf_5_25_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18443_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_145_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09944_ _10348_/A vssd1 vssd1 vccd1 vccd1 _10307_/S sky130_fd_sc_hd__buf_4
XFILLER_217_1350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_213_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09875_ _09875_/A _09875_/B vssd1 vssd1 vccd1 vccd1 _09901_/A sky130_fd_sc_hd__xnor2_2
XTAP_4007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_219_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_13 _09160_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_24 _09243_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_213_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_35 _12121_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_46 _10483_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_57 _17661_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_68 _13522_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_227_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_79 _13591_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_214_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10650_ _12966_/A _10650_/B vssd1 vssd1 vccd1 vccd1 _10779_/A sky130_fd_sc_hd__xnor2_4
XFILLER_139_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_224_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09309_ _09309_/A _10575_/A _09309_/C _09309_/D vssd1 vssd1 vccd1 vccd1 _09320_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_16_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10581_ _09344_/B _09354_/C _10391_/A _10389_/A _10036_/A _10102_/S vssd1 vssd1 vccd1
+ vccd1 _10581_/X sky130_fd_sc_hd__mux4_1
XFILLER_220_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12320_ _13210_/A vssd1 vssd1 vccd1 vccd1 _13153_/A sky130_fd_sc_hd__buf_8
XFILLER_127_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_209_wb_clk_i _17803_/CLK vssd1 vssd1 vccd1 vccd1 _18960_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_103_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_214_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12251_ _12251_/A _12285_/A _12258_/C vssd1 vssd1 vccd1 vccd1 _12251_/X sky130_fd_sc_hd__and3_1
XFILLER_5_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11202_ _11210_/A _11202_/B _11202_/C vssd1 vssd1 vccd1 vccd1 _11203_/A sky130_fd_sc_hd__and3_1
XFILLER_181_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12182_ _12180_/Y _12181_/X _12163_/X vssd1 vssd1 vccd1 vccd1 _17848_/D sky130_fd_sc_hd__o21a_1
XFILLER_79_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_218_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_190_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11133_ _11392_/B vssd1 vssd1 vccd1 vccd1 _11595_/A sky130_fd_sc_hd__clkbuf_2
X_16990_ _17078_/A vssd1 vssd1 vccd1 vccd1 _17005_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_1_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15941_ _18599_/Q _18563_/Q _15963_/S vssd1 vssd1 vccd1 vccd1 _15941_/X sky130_fd_sc_hd__mux2_1
XTAP_5220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11064_ _11064_/A vssd1 vssd1 vccd1 vccd1 _17787_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_89_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10015_ _09143_/C _09148_/B _10019_/S vssd1 vssd1 vccd1 vccd1 _10015_/X sky130_fd_sc_hd__mux2_1
XFILLER_48_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_231_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18660_ _18696_/CLK _18660_/D vssd1 vssd1 vccd1 vccd1 _18660_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_7_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15872_ _18583_/Q _18547_/Q _15879_/S vssd1 vssd1 vccd1 vccd1 _15872_/X sky130_fd_sc_hd__mux2_1
XTAP_4530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_218_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17611_ _17611_/A vssd1 vssd1 vccd1 vccd1 _18964_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14823_ _14872_/A _14827_/B vssd1 vssd1 vccd1 vccd1 _14823_/Y sky130_fd_sc_hd__nand2_1
XFILLER_40_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18591_ _18593_/CLK _18591_/D vssd1 vssd1 vccd1 vccd1 _18591_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_1208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_224_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17542_ _17544_/B _17540_/X _17541_/Y _11816_/X vssd1 vssd1 vccd1 vccd1 _18949_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_151_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14754_ _14753_/B _14752_/X _14753_/Y _14738_/X vssd1 vssd1 vccd1 vccd1 _18278_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_63_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11966_ _12028_/A _13684_/A vssd1 vssd1 vccd1 vccd1 _13434_/B sky130_fd_sc_hd__or2b_1
XTAP_3884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13705_ _13705_/A vssd1 vssd1 vccd1 vccd1 _14124_/A sky130_fd_sc_hd__buf_6
X_10917_ _10915_/X _10916_/X _10923_/S vssd1 vssd1 vccd1 vccd1 _10917_/X sky130_fd_sc_hd__mux2_1
XFILLER_17_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14685_ _17687_/A _14685_/B vssd1 vssd1 vccd1 vccd1 _16959_/A sky130_fd_sc_hd__or2_4
X_17473_ _17493_/A _17473_/B _17516_/C vssd1 vssd1 vccd1 vccd1 _17473_/X sky130_fd_sc_hd__or3_1
XFILLER_229_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11897_ _17838_/Q _12972_/A vssd1 vssd1 vccd1 vccd1 _11897_/X sky130_fd_sc_hd__and2_1
XFILLER_60_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_204_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_220_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19212_ _19212_/A _08964_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[12] sky130_fd_sc_hd__ebufn_8
X_16424_ _16473_/A vssd1 vssd1 vccd1 vccd1 _16449_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_189_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13636_ _13710_/C _13648_/B vssd1 vssd1 vccd1 vccd1 _13637_/B sky130_fd_sc_hd__or2_1
X_10848_ _10910_/C _10733_/X _10839_/X _10847_/X vssd1 vssd1 vccd1 vccd1 _10848_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_125_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19143_ _19143_/A _09052_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[13] sky130_fd_sc_hd__ebufn_8
X_16355_ _16353_/B _16352_/X _16353_/Y _16354_/X vssd1 vssd1 vccd1 vccd1 _18659_/D
+ sky130_fd_sc_hd__o211a_1
X_13567_ _13877_/A vssd1 vssd1 vccd1 vccd1 _13568_/A sky130_fd_sc_hd__buf_4
XFILLER_160_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10779_ _10779_/A vssd1 vssd1 vccd1 vccd1 _10779_/X sky130_fd_sc_hd__buf_2
XFILLER_9_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15306_ _15915_/A _15451_/C vssd1 vssd1 vccd1 vccd1 _15325_/B sky130_fd_sc_hd__nor2_1
XFILLER_201_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12518_ _12518_/A vssd1 vssd1 vccd1 vccd1 _17914_/D sky130_fd_sc_hd__clkbuf_1
X_16286_ _16285_/B _16282_/X _16285_/Y _16274_/X vssd1 vssd1 vccd1 vccd1 _18641_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_173_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13498_ _13626_/A vssd1 vssd1 vccd1 vccd1 _13592_/A sky130_fd_sc_hd__buf_8
XFILLER_121_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18025_ _18094_/CLK _18025_/D vssd1 vssd1 vccd1 vccd1 _18025_/Q sky130_fd_sc_hd__dfxtp_1
X_15237_ _15239_/B _15235_/X _15236_/Y _15224_/X vssd1 vssd1 vccd1 vccd1 _18397_/D
+ sky130_fd_sc_hd__o211a_1
X_12449_ _17903_/Q _12486_/B vssd1 vssd1 vccd1 vccd1 _12458_/A sky130_fd_sc_hd__nand2_1
XFILLER_126_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15168_ _18416_/Q _18380_/Q _15177_/S vssd1 vssd1 vccd1 vccd1 _15168_/X sky130_fd_sc_hd__mux2_1
XFILLER_160_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_113_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14119_ _18923_/Q _14017_/X _14115_/X _14118_/X vssd1 vssd1 vccd1 vccd1 _14119_/X
+ sky130_fd_sc_hd__a211o_1
X_15099_ _15107_/B _15097_/X _15098_/X _15083_/X vssd1 vssd1 vccd1 vccd1 _18363_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_141_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18927_ _18927_/CLK _18927_/D vssd1 vssd1 vccd1 vccd1 _18927_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_140_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09660_ _17975_/Q vssd1 vssd1 vccd1 vccd1 _10623_/A sky130_fd_sc_hd__clkbuf_2
X_18858_ _18858_/CLK _18858_/D vssd1 vssd1 vccd1 vccd1 _18858_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_132_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_228_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17809_ _18989_/CLK _17809_/D vssd1 vssd1 vccd1 vccd1 _17809_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_209_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09591_ _09598_/S _09591_/B vssd1 vssd1 vccd1 vccd1 _09593_/B sky130_fd_sc_hd__and2_1
XFILLER_167_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18789_ _18823_/CLK _18789_/D vssd1 vssd1 vccd1 vccd1 _18789_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_227_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_224_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XINSDIODE2_150 _18960_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_168_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_161 _18359_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_223_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_172 _18853_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_183 _09034_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_194 _09148_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_195_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_206_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_148_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09025_ _09028_/A vssd1 vssd1 vccd1 vccd1 _09025_/Y sky130_fd_sc_hd__inv_2
XFILLER_108_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_117_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_176_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09927_ _09408_/A _09408_/B _09413_/C _09418_/B _09923_/X _12123_/A vssd1 vssd1 vccd1
+ vccd1 _09927_/X sky130_fd_sc_hd__mux4_1
XFILLER_132_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09858_ _09858_/A _09858_/B vssd1 vssd1 vccd1 vccd1 _09879_/B sky130_fd_sc_hd__xor2_4
XTAP_590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09789_ _09891_/B _09891_/A vssd1 vssd1 vccd1 vccd1 _09789_/X sky130_fd_sc_hd__or2b_1
XTAP_3136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11820_ _11820_/A _11820_/B vssd1 vssd1 vccd1 vccd1 _11820_/X sky130_fd_sc_hd__and2_1
XTAP_3158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_164_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11751_ _11749_/A _11749_/C _11749_/B vssd1 vssd1 vccd1 vccd1 _11856_/C sky130_fd_sc_hd__o21a_1
XTAP_1734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_214_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10702_ _10702_/A vssd1 vssd1 vccd1 vccd1 _10856_/S sky130_fd_sc_hd__buf_4
XFILLER_14_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14470_ _14470_/A _14470_/B _14470_/C vssd1 vssd1 vccd1 vccd1 _14471_/C sky130_fd_sc_hd__nand3_1
XTAP_1778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11682_ _11503_/A _11720_/B _11593_/B _11659_/D _11681_/X vssd1 vssd1 vccd1 vccd1
+ _11683_/C sky130_fd_sc_hd__o32a_1
XFILLER_42_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_187_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_144_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13421_ _13421_/A _13648_/A vssd1 vssd1 vccd1 vccd1 _13442_/B sky130_fd_sc_hd__nand2_4
X_10633_ _10801_/S vssd1 vssd1 vccd1 vccd1 _10838_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_186_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_224_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16140_ _16147_/B _16136_/X _16138_/X _16139_/X vssd1 vssd1 vccd1 vccd1 _18609_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_220_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13352_ _09580_/A _13344_/X _11023_/X _11045_/X vssd1 vssd1 vccd1 vccd1 _18103_/D
+ sky130_fd_sc_hd__o211a_1
X_10564_ _10899_/A _10563_/X _10513_/A vssd1 vssd1 vccd1 vccd1 _10564_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_127_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12303_ _17879_/Q _11346_/A _12300_/B vssd1 vssd1 vccd1 vccd1 _12327_/B sky130_fd_sc_hd__o21a_1
X_16071_ _18630_/Q _18594_/Q _16091_/S vssd1 vssd1 vccd1 vccd1 _16071_/X sky130_fd_sc_hd__mux2_1
X_13283_ _18062_/Q _18036_/Q _18037_/Q _18039_/Q vssd1 vssd1 vccd1 vccd1 _13286_/B
+ sky130_fd_sc_hd__or4_1
X_10495_ _09093_/C _09098_/B _10495_/S vssd1 vssd1 vccd1 vccd1 _10496_/B sky130_fd_sc_hd__mux2_2
XFILLER_68_1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15022_ _15058_/A _15025_/B vssd1 vssd1 vccd1 vccd1 _15022_/Y sky130_fd_sc_hd__nand2_1
XFILLER_182_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12234_ _11896_/X _12235_/A _12228_/Y _12232_/X _12233_/X vssd1 vssd1 vccd1 vccd1
+ _17857_/D sky130_fd_sc_hd__a41o_1
XFILLER_114_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_194_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12165_ _13458_/A _12171_/C vssd1 vssd1 vccd1 vccd1 _12165_/Y sky130_fd_sc_hd__nor2_1
XFILLER_29_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11116_ _11307_/B vssd1 vssd1 vccd1 vccd1 _11452_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_1_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16973_ _16972_/B _16970_/X _16972_/Y _16964_/X vssd1 vssd1 vccd1 vccd1 _18806_/D
+ sky130_fd_sc_hd__o211a_1
X_12096_ _12982_/A _12096_/B vssd1 vssd1 vccd1 vccd1 _12097_/B sky130_fd_sc_hd__xnor2_4
XFILLER_49_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_231_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18712_ _18719_/CLK _18712_/D vssd1 vssd1 vccd1 vccd1 _18712_/Q sky130_fd_sc_hd__dfxtp_4
X_15924_ _15938_/A _15928_/B vssd1 vssd1 vccd1 vccd1 _15924_/Y sky130_fd_sc_hd__nand2_1
XTAP_5050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11047_ _17998_/Q vssd1 vssd1 vccd1 vccd1 _13394_/D sky130_fd_sc_hd__clkbuf_2
XTAP_5061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_231_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18643_ _18668_/CLK _18643_/D vssd1 vssd1 vccd1 vccd1 _18643_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_209_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15855_ _16005_/A _15892_/B vssd1 vssd1 vccd1 vccd1 _15865_/B sky130_fd_sc_hd__nor2_2
XFILLER_188_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14806_ _14928_/A vssd1 vssd1 vccd1 vccd1 _14856_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_36_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18574_ _18577_/CLK _18574_/D vssd1 vssd1 vccd1 vccd1 _18574_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_188_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15786_ _15931_/A _15844_/B vssd1 vssd1 vccd1 vccd1 _15795_/B sky130_fd_sc_hd__nor2_2
XTAP_3670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12998_ _12998_/A vssd1 vssd1 vccd1 vccd1 _17979_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_5_13_0_wb_clk_i clkbuf_4_6_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18176_/CLK
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_75_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17525_ _17524_/B _17523_/X _17524_/Y _17517_/X vssd1 vssd1 vccd1 vccd1 _18944_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_205_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14737_ _14750_/A _14742_/B vssd1 vssd1 vccd1 vccd1 _14737_/Y sky130_fd_sc_hd__nand2_1
XFILLER_166_1363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11949_ _12025_/B _11946_/X _11948_/X vssd1 vssd1 vccd1 vccd1 _12049_/A sky130_fd_sc_hd__a21o_2
XFILLER_220_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17456_ _17456_/A _17456_/B vssd1 vssd1 vccd1 vccd1 _17456_/Y sky130_fd_sc_hd__nand2_1
X_14668_ _14668_/A vssd1 vssd1 vccd1 vccd1 _14668_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_177_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16407_ _16450_/A _16407_/B vssd1 vssd1 vccd1 vccd1 _16407_/Y sky130_fd_sc_hd__nand2_1
XFILLER_203_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13619_ _13619_/A vssd1 vssd1 vccd1 vccd1 _13619_/X sky130_fd_sc_hd__buf_6
XFILLER_20_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17387_ _17448_/A vssd1 vssd1 vccd1 vccd1 _17437_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_14599_ _14687_/A vssd1 vssd1 vccd1 vccd1 _14665_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_125_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_203_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16338_ _16389_/A _16342_/B vssd1 vssd1 vccd1 vccd1 _16338_/Y sky130_fd_sc_hd__nand2_1
XFILLER_118_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_199_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16269_ _16268_/B _16267_/X _16268_/Y _16252_/X vssd1 vssd1 vccd1 vccd1 _18638_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_12_1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18008_ _18213_/CLK _18008_/D vssd1 vssd1 vccd1 vccd1 _18008_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_173_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_206_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09712_ _18251_/Q _18250_/Q _18249_/Q vssd1 vssd1 vccd1 vccd1 _09712_/X sky130_fd_sc_hd__or3_4
XFILLER_19_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_228_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_142_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_228_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09643_ _10204_/A vssd1 vssd1 vccd1 vccd1 _13353_/A sky130_fd_sc_hd__buf_2
XFILLER_132_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_215_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09574_ _09598_/S _09592_/B _09573_/X vssd1 vssd1 vccd1 vccd1 _09725_/A sky130_fd_sc_hd__a21o_1
XFILLER_167_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_215_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_93_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_212_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_93_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_223_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_221_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_221_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_1207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09008_ _09010_/A vssd1 vssd1 vccd1 vccd1 _09008_/Y sky130_fd_sc_hd__inv_2
XFILLER_3_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10280_ _09895_/X _10277_/X _10278_/X _10279_/X vssd1 vssd1 vccd1 vccd1 _10281_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_219_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13970_ _12042_/A _13962_/X _13969_/X _12028_/D vssd1 vssd1 vccd1 vccd1 _14009_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_4_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12921_ _12921_/A _12921_/B _12921_/C vssd1 vssd1 vccd1 vccd1 _12956_/A sky130_fd_sc_hd__and3_1
XFILLER_19_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15640_ _15720_/A vssd1 vssd1 vccd1 vccd1 _15640_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_46_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12852_ _12857_/C _12852_/B _12915_/B vssd1 vssd1 vccd1 vccd1 _12853_/A sky130_fd_sc_hd__and3b_1
XTAP_2221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11803_ _17790_/Q _17789_/Q _11942_/A vssd1 vssd1 vccd1 vccd1 _11976_/B sky130_fd_sc_hd__or3_1
XTAP_2254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15571_ _15570_/B _15569_/X _15570_/Y _15555_/X vssd1 vssd1 vccd1 vccd1 _18473_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_1520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12783_ _12783_/A vssd1 vssd1 vccd1 vccd1 _13066_/C sky130_fd_sc_hd__clkbuf_2
XTAP_2265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17310_ _18925_/Q _18889_/Q _17317_/S vssd1 vssd1 vccd1 vccd1 _17310_/X sky130_fd_sc_hd__mux2_1
XFILLER_14_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11734_ _11735_/A _11748_/C vssd1 vssd1 vccd1 vccd1 _11740_/A sky130_fd_sc_hd__nand2_1
XTAP_2298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14522_ _14593_/A _14620_/A vssd1 vssd1 vccd1 vccd1 _14702_/A sky130_fd_sc_hd__or2_4
XFILLER_109_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18290_ _18290_/CLK _18290_/D vssd1 vssd1 vccd1 vccd1 _18290_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_15_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_224_wb_clk_i _17803_/CLK vssd1 vssd1 vccd1 vccd1 _18989_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_1564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17241_ _17304_/A vssd1 vssd1 vccd1 vccd1 _17241_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_109_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11665_ _11669_/A _11665_/B vssd1 vssd1 vccd1 vccd1 _11848_/B sky130_fd_sc_hd__or2_1
X_14453_ _14422_/X _09505_/B _14423_/X vssd1 vssd1 vccd1 vccd1 _14453_/X sky130_fd_sc_hd__a21o_1
XFILLER_122_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_128_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13404_ _18128_/Q _13337_/A _13368_/Y vssd1 vssd1 vccd1 vccd1 _13405_/C sky130_fd_sc_hd__a21o_1
X_10616_ _10616_/A _12099_/A vssd1 vssd1 vccd1 vccd1 _10616_/Y sky130_fd_sc_hd__nor2_8
XFILLER_167_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14384_ _14384_/A _14384_/B vssd1 vssd1 vccd1 vccd1 _14399_/A sky130_fd_sc_hd__nand2_1
X_17172_ _18891_/Q _18855_/Q _17172_/S vssd1 vssd1 vccd1 vccd1 _17172_/X sky130_fd_sc_hd__mux2_1
XFILLER_155_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11596_ _11364_/A _11305_/X _11593_/Y _11595_/Y _11681_/D vssd1 vssd1 vccd1 vccd1
+ _11597_/C sky130_fd_sc_hd__o32a_1
XFILLER_183_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16123_ _16132_/A _16123_/B vssd1 vssd1 vccd1 vccd1 _16123_/Y sky130_fd_sc_hd__nand2_1
X_13335_ _18095_/Q _13313_/X _13333_/Y _13334_/X vssd1 vssd1 vccd1 vccd1 _18095_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_122_1277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10547_ _10547_/A _10547_/B _10939_/C _10547_/D vssd1 vssd1 vccd1 vccd1 _10547_/X
+ sky130_fd_sc_hd__and4_1
XFILLER_143_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16054_ _16127_/A vssd1 vssd1 vccd1 vccd1 _16208_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_143_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13266_ _13266_/A _18087_/Q vssd1 vssd1 vccd1 vccd1 _13267_/A sky130_fd_sc_hd__and2_1
X_10478_ _09270_/B _09260_/B _09260_/D _10317_/A _10462_/X _10450_/S vssd1 vssd1 vccd1
+ vccd1 _10478_/X sky130_fd_sc_hd__mux4_1
XFILLER_68_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15005_ _18339_/Q _15012_/B _15002_/X _15004_/X vssd1 vssd1 vccd1 vccd1 _18339_/D
+ sky130_fd_sc_hd__o211a_1
X_12217_ _12217_/A vssd1 vssd1 vccd1 vccd1 _17747_/A sky130_fd_sc_hd__buf_12
X_13197_ _13197_/A _18056_/Q vssd1 vssd1 vccd1 vccd1 _13198_/A sky130_fd_sc_hd__and2_1
XFILLER_9_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_69_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12148_ _17839_/Q _12171_/B _12180_/B _12146_/X _12147_/X vssd1 vssd1 vccd1 vccd1
+ _17839_/D sky130_fd_sc_hd__o2111a_1
XFILLER_2_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16956_ _18839_/Q _18803_/Q _16970_/S vssd1 vssd1 vccd1 vccd1 _16956_/X sky130_fd_sc_hd__mux2_1
X_12079_ _12079_/A vssd1 vssd1 vccd1 vccd1 _12079_/Y sky130_fd_sc_hd__inv_2
XFILLER_133_1351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15907_ _15975_/A vssd1 vssd1 vccd1 vccd1 _16041_/B sky130_fd_sc_hd__buf_2
XFILLER_37_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16887_ _17480_/A _16906_/B vssd1 vssd1 vccd1 vccd1 _16903_/B sky130_fd_sc_hd__nor2_1
XFILLER_38_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18626_ _18658_/CLK _18626_/D vssd1 vssd1 vccd1 vccd1 _18626_/Q sky130_fd_sc_hd__dfxtp_2
X_15838_ _18575_/Q _18539_/Q _15838_/S vssd1 vssd1 vccd1 vccd1 _15838_/X sky130_fd_sc_hd__mux2_1
XTAP_4190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18557_ _18557_/CLK _18557_/D vssd1 vssd1 vccd1 vccd1 _18557_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_24_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15769_ _15818_/A _15769_/B vssd1 vssd1 vccd1 vccd1 _15769_/Y sky130_fd_sc_hd__nand2_1
XFILLER_75_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17508_ _18976_/Q _18940_/Q _17515_/S vssd1 vssd1 vccd1 vccd1 _17508_/X sky130_fd_sc_hd__mux2_1
X_09290_ _18515_/Q _18514_/Q _18513_/Q vssd1 vssd1 vccd1 vccd1 _09294_/A sky130_fd_sc_hd__or3_4
XFILLER_127_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18488_ _18497_/CLK _18488_/D vssd1 vssd1 vccd1 vccd1 _18488_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_127_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17439_ _18958_/Q _18922_/Q _17447_/S vssd1 vssd1 vccd1 vccd1 _17439_/X sky130_fd_sc_hd__mux2_1
XFILLER_21_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_1344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_99_wb_clk_i clkbuf_5_28_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18482_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_133_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_217_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_28_wb_clk_i clkbuf_5_7_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18927_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_138_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_173_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_214_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_1334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_229_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_229_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_228_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09626_ _18104_/Q _10629_/A vssd1 vssd1 vccd1 vccd1 _09631_/B sky130_fd_sc_hd__xor2_1
XFILLER_43_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_1283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09557_ _10038_/B _09589_/B vssd1 vssd1 vccd1 vccd1 _12065_/A sky130_fd_sc_hd__xor2_4
XFILLER_231_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_184_1271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_197_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09488_ _18992_/Q vssd1 vssd1 vccd1 vccd1 _14507_/B sky130_fd_sc_hd__buf_6
XFILLER_54_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_221_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11450_ _11582_/A _11735_/A _11788_/B _11413_/A _11496_/A vssd1 vssd1 vccd1 vccd1
+ _11451_/B sky130_fd_sc_hd__a311o_1
XFILLER_177_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_183_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10401_ _09314_/A _09319_/B _09314_/D _09314_/C _12124_/A _10291_/X vssd1 vssd1 vccd1
+ vccd1 _10401_/X sky130_fd_sc_hd__mux4_2
X_11381_ _11828_/B vssd1 vssd1 vccd1 vccd1 _11525_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_109_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_164_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13120_ _13142_/A vssd1 vssd1 vccd1 vccd1 _13129_/A sky130_fd_sc_hd__clkbuf_1
X_10332_ _09227_/A _09237_/B _10826_/A _09227_/D _09972_/B _09948_/A vssd1 vssd1 vccd1
+ vccd1 _10332_/X sky130_fd_sc_hd__mux4_1
XFILLER_11_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13051_ _18005_/Q _18004_/Q _18003_/Q vssd1 vssd1 vccd1 vccd1 _13058_/B sky130_fd_sc_hd__a21boi_1
X_10263_ _10238_/A _10238_/B _10211_/A vssd1 vssd1 vccd1 vccd1 _10264_/B sky130_fd_sc_hd__a21o_1
XFILLER_133_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12002_ _12041_/C _12026_/C _12026_/B vssd1 vssd1 vccd1 vccd1 _12021_/B sky130_fd_sc_hd__o21ai_4
XFILLER_79_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10194_ _18099_/Q _17973_/Q vssd1 vssd1 vccd1 vccd1 _10204_/B sky130_fd_sc_hd__xor2_2
XFILLER_120_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16810_ _16960_/B vssd1 vssd1 vccd1 vccd1 _16866_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_121_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17790_ _18986_/CLK _17790_/D vssd1 vssd1 vccd1 vccd1 _17790_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_19_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16741_ _16743_/B _16738_/X _16739_/Y _16740_/X vssd1 vssd1 vccd1 vccd1 _18754_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_207_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13953_ _18490_/Q _13733_/X _13949_/X _13952_/X vssd1 vssd1 vccd1 vccd1 _13953_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_19_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_207_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12904_ _17964_/Q _17965_/Q _12904_/C vssd1 vssd1 vccd1 vccd1 _12908_/B sky130_fd_sc_hd__and3_1
XFILLER_207_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16672_ _16672_/A _16796_/C vssd1 vssd1 vccd1 vccd1 _16686_/B sky130_fd_sc_hd__nor2_2
XFILLER_59_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13884_ _18964_/Q _13739_/X _13703_/A _18979_/Q vssd1 vssd1 vccd1 vccd1 _13884_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_207_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18411_ _18432_/CLK _18411_/D vssd1 vssd1 vccd1 vccd1 _18411_/Q sky130_fd_sc_hd__dfxtp_1
X_15623_ _15717_/A vssd1 vssd1 vccd1 vccd1 _15642_/S sky130_fd_sc_hd__clkbuf_2
XTAP_2040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_146_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12835_ _12835_/A _12835_/B _12835_/C _12835_/D vssd1 vssd1 vccd1 vccd1 _12835_/X
+ sky130_fd_sc_hd__or4_1
XTAP_2051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18342_ _18343_/CLK _18342_/D vssd1 vssd1 vccd1 vccd1 _18342_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_43_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15554_ _15566_/A _15558_/B vssd1 vssd1 vccd1 vccd1 _15554_/Y sky130_fd_sc_hd__nand2_1
XFILLER_163_1322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_187_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12766_ _12718_/X _12762_/X _12765_/Y vssd1 vssd1 vccd1 vccd1 _17940_/D sky130_fd_sc_hd__a21oi_1
XFILLER_61_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_187_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14505_ _14505_/A vssd1 vssd1 vccd1 vccd1 _18226_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18273_ _18299_/CLK _18273_/D vssd1 vssd1 vccd1 vccd1 _18273_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11717_ _11820_/A _11860_/A vssd1 vssd1 vccd1 vccd1 _11717_/Y sky130_fd_sc_hd__nor2_1
X_15485_ _15487_/B _15483_/X _15484_/Y _15474_/X vssd1 vssd1 vccd1 vccd1 _18451_/D
+ sky130_fd_sc_hd__o211a_1
X_12697_ _17939_/Q _12697_/B vssd1 vssd1 vccd1 vccd1 _12707_/B sky130_fd_sc_hd__nor2_1
XFILLER_204_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17224_ _17273_/A _17230_/B vssd1 vssd1 vccd1 vccd1 _17224_/Y sky130_fd_sc_hd__nand2_1
X_11648_ _11671_/B vssd1 vssd1 vccd1 vccd1 _11648_/X sky130_fd_sc_hd__clkbuf_2
X_14436_ _14436_/A vssd1 vssd1 vccd1 vccd1 _14436_/X sky130_fd_sc_hd__buf_8
XFILLER_200_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17155_ _18887_/Q _18851_/Q _17172_/S vssd1 vssd1 vccd1 vccd1 _17155_/X sky130_fd_sc_hd__mux2_1
XFILLER_190_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11579_ _11844_/A _11564_/X _11574_/X _11578_/Y vssd1 vssd1 vccd1 vccd1 _11579_/X
+ sky130_fd_sc_hd__a211o_1
X_14367_ _14373_/A _14381_/A _18185_/Q vssd1 vssd1 vccd1 vccd1 _14367_/X sky130_fd_sc_hd__or3b_1
XFILLER_196_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16106_ _16130_/A _16109_/B vssd1 vssd1 vccd1 vccd1 _16106_/Y sky130_fd_sc_hd__nand2_1
XFILLER_128_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13318_ _13318_/A _13318_/B _13318_/C vssd1 vssd1 vccd1 vccd1 _13318_/X sky130_fd_sc_hd__or3_1
X_17086_ _17091_/B _17083_/X _17085_/X _17076_/X vssd1 vssd1 vccd1 vccd1 _18834_/D
+ sky130_fd_sc_hd__o211a_1
X_14298_ _14294_/X _14296_/Y _14349_/A vssd1 vssd1 vccd1 vccd1 _14298_/X sky130_fd_sc_hd__mux2_1
XFILLER_170_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16037_ _16039_/B _16035_/X _16036_/Y _16028_/X vssd1 vssd1 vccd1 vccd1 _18586_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_171_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13249_ _13255_/A _18079_/Q vssd1 vssd1 vccd1 vccd1 _13250_/A sky130_fd_sc_hd__and2_1
XFILLER_42_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17988_ _18044_/CLK _17988_/D vssd1 vssd1 vccd1 vccd1 _17988_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_96_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_211_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16939_ _16954_/A _16943_/B vssd1 vssd1 vccd1 vccd1 _16939_/Y sky130_fd_sc_hd__nand2_1
XFILLER_38_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_226_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_146_wb_clk_i clkbuf_5_26_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18308_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_38_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09411_ _18332_/Q _18331_/Q _18330_/Q vssd1 vssd1 vccd1 vccd1 _09413_/C sky130_fd_sc_hd__or3_2
X_18609_ _18633_/CLK _18609_/D vssd1 vssd1 vccd1 vccd1 _18609_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_16_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09342_ _18446_/Q _18445_/Q _18444_/Q vssd1 vssd1 vccd1 vccd1 _09344_/C sky130_fd_sc_hd__or3_2
XFILLER_179_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_221_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09273_ _18860_/Q _18859_/Q _18858_/Q vssd1 vssd1 vccd1 vccd1 _09277_/A sky130_fd_sc_hd__or3_2
XFILLER_194_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_194_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_1283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_1351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_5_6_0_wb_clk_i clkbuf_5_7_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_5_6_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_107_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19115__86 vssd1 vssd1 vccd1 vccd1 _19115__86/HI _19223_/A sky130_fd_sc_hd__conb_1
XFILLER_162_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_1278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08988_ _08991_/A vssd1 vssd1 vccd1 vccd1 _08988_/Y sky130_fd_sc_hd__inv_2
XTAP_4926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_1330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_228_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10950_ _09952_/A _09402_/B _09397_/A _09392_/D _09689_/X _10942_/A vssd1 vssd1 vccd1
+ vccd1 _10950_/X sky130_fd_sc_hd__mux4_1
XFILLER_216_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09609_ _09609_/A _09609_/B vssd1 vssd1 vccd1 vccd1 _09610_/B sky130_fd_sc_hd__xnor2_2
X_10881_ _09365_/B _09370_/C _09365_/D _09360_/D _10851_/A _10852_/A vssd1 vssd1 vccd1
+ vccd1 _10881_/X sky130_fd_sc_hd__mux4_1
XFILLER_83_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12620_ _12619_/A _12619_/B _12569_/A vssd1 vssd1 vccd1 vccd1 _12620_/Y sky130_fd_sc_hd__a21oi_1
XPHY_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_189_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12551_ _12564_/A vssd1 vssd1 vccd1 vccd1 _12588_/B sky130_fd_sc_hd__clkbuf_2
XPHY_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_196_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11502_ _11491_/A _11371_/X _11394_/X _11493_/X _11501_/X vssd1 vssd1 vccd1 vccd1
+ _11502_/X sky130_fd_sc_hd__o311a_1
XFILLER_157_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15270_ _15270_/A vssd1 vssd1 vccd1 vccd1 _15285_/S sky130_fd_sc_hd__clkbuf_2
X_12482_ _12480_/Y _12484_/B _12490_/A vssd1 vssd1 vccd1 vccd1 _12482_/X sky130_fd_sc_hd__o21a_1
XFILLER_40_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11433_ _11423_/A _12323_/A _19029_/Q vssd1 vssd1 vccd1 vccd1 _11433_/X sky130_fd_sc_hd__and3b_1
X_14221_ _14323_/B vssd1 vssd1 vccd1 vccd1 _14305_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_172_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14152_ _13637_/Y _14128_/X _14151_/X vssd1 vssd1 vccd1 vccd1 _14152_/X sky130_fd_sc_hd__a21o_1
X_11364_ _11364_/A _11364_/B vssd1 vssd1 vccd1 vccd1 _11468_/B sky130_fd_sc_hd__nor2_1
XFILLER_138_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_193_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_217_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13103_ _13107_/A _18013_/Q vssd1 vssd1 vccd1 vccd1 _13104_/A sky130_fd_sc_hd__and2_1
X_10315_ _09260_/A _09270_/C _09270_/D _09265_/D _10291_/X _09935_/X vssd1 vssd1 vccd1
+ vccd1 _10315_/X sky130_fd_sc_hd__mux4_1
X_14083_ _18467_/Q _13525_/A _13621_/X _18470_/Q vssd1 vssd1 vccd1 vccd1 _14083_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_152_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18960_ _18960_/CLK _18960_/D vssd1 vssd1 vccd1 vccd1 _18960_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_98_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11295_ _11336_/A _11336_/B _11333_/A vssd1 vssd1 vccd1 vccd1 _11312_/B sky130_fd_sc_hd__nand3_1
XFILLER_4_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17911_ _17911_/CLK _17911_/D vssd1 vssd1 vccd1 vccd1 _17911_/Q sky130_fd_sc_hd__dfxtp_1
X_13034_ _13016_/X _13000_/A _12935_/X _13210_/A vssd1 vssd1 vccd1 vccd1 _13034_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_152_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10246_ _10246_/A _10246_/B vssd1 vssd1 vccd1 vccd1 _11910_/A sky130_fd_sc_hd__or2_1
XFILLER_117_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18891_ _18893_/CLK _18891_/D vssd1 vssd1 vccd1 vccd1 _18891_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_133_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17842_ _17890_/CLK _17842_/D vssd1 vssd1 vccd1 vccd1 _17842_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_65_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10177_ _10175_/A _10175_/B _10147_/A vssd1 vssd1 vccd1 vccd1 _10179_/A sky130_fd_sc_hd__a21oi_2
XFILLER_78_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17773_ _19031_/Q _12284_/X _14436_/X vssd1 vssd1 vccd1 vccd1 _19031_/D sky130_fd_sc_hd__o21a_1
X_14985_ _15277_/A _14985_/B vssd1 vssd1 vccd1 vccd1 _14995_/B sky130_fd_sc_hd__nor2_2
XFILLER_208_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16724_ _16760_/A vssd1 vssd1 vccd1 vccd1 _16724_/X sky130_fd_sc_hd__clkbuf_2
X_13936_ _18334_/Q _13738_/X _13934_/X _13935_/X vssd1 vssd1 vccd1 vccd1 _13936_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_130_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_219_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_228_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_223_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_207_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16655_ _16695_/A _16658_/B vssd1 vssd1 vccd1 vccd1 _16655_/Y sky130_fd_sc_hd__nand2_1
XFILLER_34_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13867_ _12027_/B _13855_/X _13866_/X _13434_/C vssd1 vssd1 vccd1 vccd1 _13867_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_179_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15606_ _15605_/B _15604_/X _15605_/Y _15595_/X vssd1 vssd1 vccd1 vccd1 _18482_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_16_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12818_ _12533_/Y _17946_/Q _17963_/Q _12662_/A _12817_/Y vssd1 vssd1 vccd1 vccd1
+ _12818_/X sky130_fd_sc_hd__a221o_1
X_16586_ _18715_/Q _16589_/B _16585_/Y _16581_/X vssd1 vssd1 vccd1 vccd1 _18715_/D
+ sky130_fd_sc_hd__o211a_1
X_13798_ _18351_/Q _13781_/A _13721_/A _18366_/Q vssd1 vssd1 vccd1 vccd1 _13798_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_37_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18325_ _18350_/CLK _18325_/D vssd1 vssd1 vccd1 vccd1 _18325_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_128_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15537_ _18464_/Q _15534_/B _15534_/Y _15536_/X vssd1 vssd1 vccd1 vccd1 _18464_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_1180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_231_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12749_ _18033_/Q _18032_/Q _18035_/Q _18034_/Q vssd1 vssd1 vccd1 vccd1 _12752_/A
+ sky130_fd_sc_hd__and4_1
XTAP_1191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18256_ _18266_/CLK _18256_/D vssd1 vssd1 vccd1 vccd1 _18256_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_8_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15468_ _15597_/B vssd1 vssd1 vccd1 vccd1 _15515_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_148_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17207_ _17256_/A _17493_/B _17234_/C vssd1 vssd1 vccd1 vccd1 _17207_/X sky130_fd_sc_hd__or3_1
XFILLER_128_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14419_ _18195_/Q _14418_/X _14401_/X _09498_/B vssd1 vssd1 vccd1 vccd1 _14420_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_200_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18187_ _18230_/CLK _18187_/D vssd1 vssd1 vccd1 vccd1 _18187_/Q sky130_fd_sc_hd__dfxtp_1
X_15399_ _18469_/Q _18433_/Q _15412_/S vssd1 vssd1 vccd1 vccd1 _15399_/X sky130_fd_sc_hd__mux2_1
XFILLER_162_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17138_ _18883_/Q _18847_/Q _17151_/S vssd1 vssd1 vccd1 vccd1 _17138_/X sky130_fd_sc_hd__mux2_1
XFILLER_171_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17069_ _17068_/B _17067_/X _17068_/Y _17057_/X vssd1 vssd1 vccd1 vccd1 _18830_/D
+ sky130_fd_sc_hd__o211a_1
X_09960_ _09365_/A _09370_/B _10883_/A _09360_/C _10285_/S _09959_/X vssd1 vssd1 vccd1
+ vccd1 _09960_/X sky130_fd_sc_hd__mux4_1
XFILLER_104_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_98_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09891_ _09891_/A _09891_/B vssd1 vssd1 vccd1 vccd1 _09892_/B sky130_fd_sc_hd__xor2_2
XTAP_931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_214_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_226_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_214_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_226_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_214_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_213_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_198_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09325_ _18539_/Q _18538_/Q _18537_/Q vssd1 vssd1 vccd1 vccd1 _09327_/C sky130_fd_sc_hd__or3_1
XFILLER_159_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_221_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09256_ _18962_/Q _18961_/Q _18960_/Q vssd1 vssd1 vccd1 vccd1 _09260_/A sky130_fd_sc_hd__or3_2
XFILLER_194_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_43_wb_clk_i clkbuf_5_16_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18778_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_181_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09187_ _09187_/A _09187_/B _09187_/C vssd1 vssd1 vccd1 vccd1 _09187_/Y sky130_fd_sc_hd__nand3_1
XFILLER_175_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_218_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10100_ _10029_/S _10095_/X _10099_/X _10010_/A vssd1 vssd1 vccd1 vccd1 _10100_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_108_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11080_ _11970_/A vssd1 vssd1 vccd1 vccd1 _11984_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_68_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10031_ _09720_/X _10021_/X _10030_/X _10895_/A vssd1 vssd1 vccd1 vccd1 _10031_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_5424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_191_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_194_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14770_ _17473_/B _14843_/C vssd1 vssd1 vccd1 vccd1 _14777_/B sky130_fd_sc_hd__nor2_2
XTAP_4789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11982_ _12022_/A _13434_/A _13421_/A vssd1 vssd1 vccd1 vccd1 _12055_/C sky130_fd_sc_hd__or3b_4
XFILLER_29_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_216_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13721_ _13721_/A vssd1 vssd1 vccd1 vccd1 _13721_/X sky130_fd_sc_hd__buf_6
XFILLER_17_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10933_ _09304_/D _09299_/D _09294_/C _09299_/B _10495_/S _10522_/X vssd1 vssd1 vccd1
+ vccd1 _10933_/X sky130_fd_sc_hd__mux4_1
XFILLER_71_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16440_ _18680_/Q _16439_/B _16439_/Y _16437_/X vssd1 vssd1 vccd1 vccd1 _18680_/D
+ sky130_fd_sc_hd__o211a_1
X_13652_ _13652_/A vssd1 vssd1 vccd1 vccd1 _13781_/A sky130_fd_sc_hd__buf_4
X_10864_ _10864_/A vssd1 vssd1 vccd1 vccd1 _14247_/A sky130_fd_sc_hd__buf_2
XFILLER_73_1311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_220_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12603_ _12529_/X _12600_/Y _12601_/X _12602_/Y vssd1 vssd1 vccd1 vccd1 _17924_/D
+ sky130_fd_sc_hd__a31o_1
X_16371_ _16371_/A _16666_/B _16422_/C vssd1 vssd1 vccd1 vccd1 _16371_/X sky130_fd_sc_hd__or3_1
XPHY_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13583_ _13583_/A vssd1 vssd1 vccd1 vccd1 _13760_/A sky130_fd_sc_hd__clkbuf_8
XPHY_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10795_ _10795_/A _10813_/B vssd1 vssd1 vccd1 vccd1 _10795_/X sky130_fd_sc_hd__or2_1
XFILLER_213_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18110_ _18110_/CLK _18110_/D vssd1 vssd1 vccd1 vccd1 _18110_/Q sky130_fd_sc_hd__dfxtp_1
X_15322_ _18452_/Q _18416_/Q _15334_/S vssd1 vssd1 vccd1 vccd1 _15322_/X sky130_fd_sc_hd__mux2_1
XPHY_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_223_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12534_ _17920_/Q _17917_/Q vssd1 vssd1 vccd1 vccd1 _12535_/B sky130_fd_sc_hd__xnor2_2
XFILLER_160_1358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_219_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18041_ _18052_/CLK _18041_/D vssd1 vssd1 vccd1 vccd1 _18041_/Q sky130_fd_sc_hd__dfxtp_1
X_15253_ _15303_/A _15253_/B vssd1 vssd1 vccd1 vccd1 _15253_/Y sky130_fd_sc_hd__nand2_1
XFILLER_8_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12465_ _12466_/B _12466_/C _12477_/C vssd1 vssd1 vccd1 vccd1 _12465_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_149_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14204_ _18996_/Q _14204_/B vssd1 vssd1 vccd1 vccd1 _14205_/A sky130_fd_sc_hd__and2b_1
XFILLER_125_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11416_ _17882_/Q vssd1 vssd1 vccd1 vccd1 _11423_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_15184_ _15184_/A _15229_/B vssd1 vssd1 vccd1 vccd1 _15195_/B sky130_fd_sc_hd__nor2_1
X_12396_ _12397_/A _12397_/B _12397_/C vssd1 vssd1 vccd1 vccd1 _12406_/B sky130_fd_sc_hd__o21a_1
X_14135_ _18302_/Q _13612_/A _14027_/A _18293_/Q _14134_/X vssd1 vssd1 vccd1 vccd1
+ _14135_/X sky130_fd_sc_hd__a221o_4
X_11347_ _11622_/A _11323_/X _11325_/Y _11342_/X _11346_/Y vssd1 vssd1 vccd1 vccd1
+ _11347_/X sky130_fd_sc_hd__o311a_1
XFILLER_193_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14066_ _13434_/A _14035_/X _14050_/X _14065_/X vssd1 vssd1 vccd1 vccd1 _14066_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_152_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11278_ _11970_/A _17793_/Q _11926_/B vssd1 vssd1 vccd1 vccd1 _11281_/B sky130_fd_sc_hd__or3_2
X_18943_ _18953_/CLK _18943_/D vssd1 vssd1 vccd1 vccd1 _18943_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_80_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10229_ _10559_/S vssd1 vssd1 vccd1 vccd1 _10518_/A sky130_fd_sc_hd__buf_4
X_13017_ _13016_/X _12961_/A _12718_/X _11891_/X vssd1 vssd1 vccd1 vccd1 _13017_/X
+ sky130_fd_sc_hd__a31o_1
X_18874_ _18875_/CLK _18874_/D vssd1 vssd1 vccd1 vccd1 _18874_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_79_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_228_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17825_ _18157_/CLK _17825_/D vssd1 vssd1 vccd1 vccd1 _17825_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_67_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_227_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xhold1 hold1/A vssd1 vssd1 vccd1 vccd1 hold1/X sky130_fd_sc_hd__clkdlybuf4s25_1
XTAP_5980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17756_ _17756_/A _19022_/Q vssd1 vssd1 vccd1 vccd1 _17757_/A sky130_fd_sc_hd__and2_1
XFILLER_78_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14968_ _14992_/A _14971_/B vssd1 vssd1 vccd1 vccd1 _14968_/Y sky130_fd_sc_hd__nand2_1
XFILLER_35_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16707_ _16828_/A vssd1 vssd1 vccd1 vccd1 _16752_/A sky130_fd_sc_hd__clkbuf_2
X_13919_ _18766_/Q _13940_/A _14030_/A _18763_/Q vssd1 vssd1 vccd1 vccd1 _13919_/X
+ sky130_fd_sc_hd__a22o_1
X_17687_ _17687_/A _17687_/B vssd1 vssd1 vccd1 vccd1 _17687_/Y sky130_fd_sc_hd__nor2_1
X_14899_ _18350_/Q _18314_/Q _14905_/S vssd1 vssd1 vccd1 vccd1 _14899_/X sky130_fd_sc_hd__mux2_1
XFILLER_78_1266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_223_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16638_ _16678_/A _16785_/B _16652_/C vssd1 vssd1 vccd1 vccd1 _16638_/X sky130_fd_sc_hd__or3_1
XFILLER_62_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_222_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_222_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16569_ _16575_/B _16565_/X _16568_/X _16559_/X vssd1 vssd1 vccd1 vccd1 _18711_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_22_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09110_ _18749_/Q _18748_/Q _18747_/Q vssd1 vssd1 vccd1 vccd1 _09114_/A sky130_fd_sc_hd__or3_4
XFILLER_188_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18308_ _18308_/CLK _18308_/D vssd1 vssd1 vccd1 vccd1 _18308_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_128_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09041_ _09053_/A vssd1 vssd1 vccd1 vccd1 _09046_/A sky130_fd_sc_hd__buf_12
XFILLER_191_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18239_ _18263_/CLK _18239_/D vssd1 vssd1 vccd1 vccd1 _18239_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_198_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_1321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09943_ _10333_/S vssd1 vssd1 vccd1 vccd1 _12128_/A sky130_fd_sc_hd__buf_4
XFILLER_132_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_217_1362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_225_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_225_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_161_wb_clk_i clkbuf_5_11_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18061_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_09874_ _09874_/A _09880_/A vssd1 vssd1 vccd1 vccd1 _09875_/B sky130_fd_sc_hd__xnor2_1
XTAP_761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_14 _09170_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_25 _09253_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_36 _12123_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINSDIODE2_47 _10484_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_58 _16891_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_69 _13522_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_213_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_202_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_183_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09308_ _18452_/Q _18451_/Q _18450_/Q vssd1 vssd1 vccd1 vccd1 _09309_/D sky130_fd_sc_hd__or3_4
X_10580_ _09349_/A _09354_/A _09344_/A _09349_/B _10568_/X _10025_/A vssd1 vssd1 vccd1
+ vccd1 _10580_/X sky130_fd_sc_hd__mux4_1
XFILLER_10_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_107_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09239_ _18884_/Q _18883_/Q _18882_/Q vssd1 vssd1 vccd1 vccd1 _09243_/A sky130_fd_sc_hd__or3_4
XFILLER_166_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_222_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_182_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12250_ _11639_/A _11648_/X _12251_/A vssd1 vssd1 vccd1 vccd1 _12250_/X sky130_fd_sc_hd__a21o_1
XFILLER_5_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11201_ _11201_/A _11205_/C vssd1 vssd1 vccd1 vccd1 _11202_/C sky130_fd_sc_hd__nand2_1
XFILLER_107_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12181_ _17848_/Q _12172_/B _12165_/Y vssd1 vssd1 vccd1 vccd1 _12181_/X sky130_fd_sc_hd__a21o_1
XFILLER_107_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_122_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11132_ _11453_/A vssd1 vssd1 vccd1 vccd1 _11392_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_190_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_1204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15940_ _16014_/A vssd1 vssd1 vccd1 vccd1 _15963_/S sky130_fd_sc_hd__clkbuf_2
XTAP_5210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11063_ _13427_/A _11224_/A _12272_/A vssd1 vssd1 vccd1 vccd1 _11064_/A sky130_fd_sc_hd__mux2_1
XFILLER_95_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10014_ _10096_/S vssd1 vssd1 vccd1 vccd1 _10019_/S sky130_fd_sc_hd__buf_2
XFILLER_23_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_209_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15871_ _15876_/B _15868_/X _15870_/X _15861_/X vssd1 vssd1 vccd1 vccd1 _18546_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_4520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17610_ _17610_/A _17610_/B vssd1 vssd1 vccd1 vccd1 _17611_/A sky130_fd_sc_hd__and2_1
XTAP_5298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14822_ _14944_/A vssd1 vssd1 vccd1 vccd1 _14872_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_76_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18590_ _18590_/CLK _18590_/D vssd1 vssd1 vccd1 vccd1 _18590_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_4564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17541_ _17541_/A _17544_/B vssd1 vssd1 vccd1 vccd1 _17541_/Y sky130_fd_sc_hd__nand2_1
XFILLER_205_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14753_ _14753_/A _14753_/B vssd1 vssd1 vccd1 vccd1 _14753_/Y sky130_fd_sc_hd__nand2_1
XFILLER_91_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_229_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11965_ _12007_/A _12020_/B _11960_/B vssd1 vssd1 vccd1 vccd1 _13684_/A sky130_fd_sc_hd__or3b_2
XTAP_3885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13704_ _18765_/Q _13940_/A _14030_/A _18762_/Q vssd1 vssd1 vccd1 vccd1 _13704_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_204_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10916_ _09314_/C _09314_/D _09319_/B _09314_/A _10518_/X _10236_/A vssd1 vssd1 vccd1
+ vccd1 _10916_/X sky130_fd_sc_hd__mux4_1
XFILLER_44_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17472_ _17472_/A vssd1 vssd1 vccd1 vccd1 _17516_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_14684_ _18263_/Q _14683_/B _14683_/Y _14668_/X vssd1 vssd1 vccd1 vccd1 _18263_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_225_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_205_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11896_ _14457_/B vssd1 vssd1 vccd1 vccd1 _11896_/X sky130_fd_sc_hd__buf_8
XFILLER_189_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19211_ _19211_/A _08963_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[11] sky130_fd_sc_hd__ebufn_8
XFILLER_32_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16423_ _16429_/B _16421_/X _16422_/X _16418_/X vssd1 vssd1 vccd1 vccd1 _18675_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_204_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13635_ _13635_/A _13693_/A vssd1 vssd1 vccd1 vccd1 _13648_/B sky130_fd_sc_hd__or2b_1
X_10847_ _10679_/A _10840_/X _10844_/X _10846_/X vssd1 vssd1 vccd1 vccd1 _10847_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_38_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_1280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19142_ _19142_/A _09054_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[12] sky130_fd_sc_hd__ebufn_8
XFILLER_73_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16354_ _16354_/A vssd1 vssd1 vccd1 vccd1 _16354_/X sky130_fd_sc_hd__clkbuf_2
X_13566_ _13566_/A vssd1 vssd1 vccd1 vccd1 _13877_/A sky130_fd_sc_hd__buf_6
X_10778_ _10818_/A _10775_/X _10777_/X _10805_/B vssd1 vssd1 vccd1 vccd1 _10778_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_34_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15305_ _16823_/A vssd1 vssd1 vccd1 vccd1 _15915_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_199_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12517_ _12517_/A _12517_/B vssd1 vssd1 vccd1 vccd1 _12518_/A sky130_fd_sc_hd__and2_1
X_16285_ _16329_/A _16285_/B vssd1 vssd1 vccd1 vccd1 _16285_/Y sky130_fd_sc_hd__nand2_1
XFILLER_200_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13497_ _13763_/A vssd1 vssd1 vccd1 vccd1 _13626_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_201_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18024_ _18030_/CLK _18024_/D vssd1 vssd1 vccd1 vccd1 _18024_/Q sky130_fd_sc_hd__dfxtp_1
X_15236_ _15236_/A _15239_/B vssd1 vssd1 vccd1 vccd1 _15236_/Y sky130_fd_sc_hd__nand2_1
XFILLER_172_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12448_ _12443_/Y _12452_/B _12447_/X _12472_/A vssd1 vssd1 vccd1 vccd1 _17902_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_201_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_201_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15167_ _15169_/B _15164_/X _15165_/Y _15166_/X vssd1 vssd1 vccd1 vccd1 _18379_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_160_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12379_ _12459_/A _12379_/B _12379_/C vssd1 vssd1 vccd1 vccd1 _12380_/A sky130_fd_sc_hd__and3_1
XFILLER_158_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14118_ _18935_/Q _13525_/X _14116_/X _14117_/X vssd1 vssd1 vccd1 vccd1 _14118_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_10_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15098_ _15098_/A _15243_/B _15112_/C vssd1 vssd1 vccd1 vccd1 _15098_/X sky130_fd_sc_hd__or3_1
XFILLER_114_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14049_ _18554_/Q _14015_/A _14043_/X _14048_/X vssd1 vssd1 vccd1 vccd1 _14049_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_140_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18926_ _18926_/CLK _18926_/D vssd1 vssd1 vccd1 vccd1 _18926_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_80_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18857_ _18862_/CLK _18857_/D vssd1 vssd1 vccd1 vccd1 _18857_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_228_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_227_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17808_ _18191_/CLK _17808_/D vssd1 vssd1 vccd1 vccd1 _17808_/Q sky130_fd_sc_hd__dfxtp_1
X_09590_ _09555_/B _09590_/B vssd1 vssd1 vccd1 vccd1 _09593_/A sky130_fd_sc_hd__and2b_1
X_18788_ _18788_/CLK _18788_/D vssd1 vssd1 vccd1 vccd1 _18788_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_95_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17739_ _17745_/A _19014_/Q vssd1 vssd1 vccd1 vccd1 _17740_/A sky130_fd_sc_hd__and2_1
XFILLER_78_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_224_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XINSDIODE2_140 _15921_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_151 _18419_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINSDIODE2_162 _18359_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_168_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XINSDIODE2_173 _18743_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_223_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XINSDIODE2_184 _09098_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_195 _09153_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_176_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_164_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09024_ _09028_/A vssd1 vssd1 vccd1 vccd1 _09024_/Y sky130_fd_sc_hd__inv_2
XFILLER_163_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_172_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09926_ _12124_/A vssd1 vssd1 vccd1 vccd1 _12123_/A sky130_fd_sc_hd__buf_6
XFILLER_98_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09857_ _09822_/A _09846_/B _09846_/A vssd1 vssd1 vccd1 vccd1 _09879_/A sky130_fd_sc_hd__a21boi_4
XTAP_591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_1368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09788_ _09805_/A _09793_/B vssd1 vssd1 vccd1 vccd1 _09891_/A sky130_fd_sc_hd__xnor2_2
XTAP_3126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11750_ _11733_/Y _11824_/A _11741_/X _11856_/A _11856_/B vssd1 vssd1 vccd1 vccd1
+ _11750_/Y sky130_fd_sc_hd__a311oi_1
XTAP_1724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10701_ _10701_/A vssd1 vssd1 vccd1 vccd1 _10702_/A sky130_fd_sc_hd__buf_4
XTAP_1757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11681_ _11497_/B _12089_/B _11681_/C _11681_/D vssd1 vssd1 vccd1 vccd1 _11681_/X
+ sky130_fd_sc_hd__and4b_1
XTAP_1779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_201_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_230_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_224_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13420_ _13420_/A vssd1 vssd1 vccd1 vccd1 _13648_/A sky130_fd_sc_hd__buf_2
XFILLER_197_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10632_ _12966_/A _10650_/B vssd1 vssd1 vccd1 vccd1 _10801_/S sky130_fd_sc_hd__xor2_4
XFILLER_220_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_224_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10563_ _10443_/A _10561_/X _10562_/X _10183_/A vssd1 vssd1 vccd1 vccd1 _10563_/X
+ sky130_fd_sc_hd__a22o_2
X_13351_ _09743_/A _13344_/X _11023_/X _11031_/X vssd1 vssd1 vccd1 vccd1 _18102_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_194_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_139_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12302_ _12299_/B _12292_/B _12301_/Y _12219_/X vssd1 vssd1 vccd1 vccd1 _17875_/D
+ sky130_fd_sc_hd__o211a_1
X_16070_ _16173_/A vssd1 vssd1 vccd1 vccd1 _16091_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_127_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10494_ _10494_/A vssd1 vssd1 vccd1 vccd1 _10495_/S sky130_fd_sc_hd__buf_2
XFILLER_5_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13282_ _18029_/Q _18028_/Q _18031_/Q _18030_/Q vssd1 vssd1 vccd1 vccd1 _13286_/A
+ sky130_fd_sc_hd__or4_1
XFILLER_136_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15021_ _18379_/Q _18343_/Q _15033_/S vssd1 vssd1 vccd1 vccd1 _15021_/X sky130_fd_sc_hd__mux2_1
XFILLER_108_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12233_ _12233_/A _12285_/A _12233_/C vssd1 vssd1 vccd1 vccd1 _12233_/X sky130_fd_sc_hd__and3_1
XFILLER_30_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12164_ _12160_/Y _12161_/X _12163_/X vssd1 vssd1 vccd1 vccd1 _17843_/D sky130_fd_sc_hd__o21a_1
XFILLER_151_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11115_ _17798_/Q vssd1 vssd1 vccd1 vccd1 _11307_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_19076__47 vssd1 vssd1 vccd1 vccd1 _19076__47/HI _19170_/A sky130_fd_sc_hd__conb_1
X_16972_ _17035_/A _16972_/B vssd1 vssd1 vccd1 vccd1 _16972_/Y sky130_fd_sc_hd__nand2_1
XFILLER_122_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12095_ _12095_/A _12095_/B _12095_/C _12095_/D vssd1 vssd1 vccd1 vccd1 _12104_/A
+ sky130_fd_sc_hd__or4_1
XFILLER_110_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_150_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15923_ _18595_/Q _18559_/Q _15937_/S vssd1 vssd1 vccd1 vccd1 _15923_/X sky130_fd_sc_hd__mux2_1
X_18711_ _18722_/CLK _18711_/D vssd1 vssd1 vccd1 vccd1 _18711_/Q sky130_fd_sc_hd__dfxtp_4
X_11046_ _17999_/Q vssd1 vssd1 vccd1 vccd1 _13375_/A sky130_fd_sc_hd__buf_2
XFILLER_231_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18642_ _18668_/CLK _18642_/D vssd1 vssd1 vccd1 vccd1 _18642_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_5084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_231_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15854_ _15853_/B _15852_/X _15853_/Y _15842_/X vssd1 vssd1 vccd1 vccd1 _18542_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_4350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_225_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_225_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14805_ _18327_/Q _18291_/Q _14809_/S vssd1 vssd1 vccd1 vccd1 _14805_/X sky130_fd_sc_hd__mux2_1
XFILLER_18_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18573_ _18577_/CLK _18573_/D vssd1 vssd1 vccd1 vccd1 _18573_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_4394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15785_ _15821_/A vssd1 vssd1 vccd1 vccd1 _15844_/B sky130_fd_sc_hd__buf_2
XTAP_3660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12997_ _13049_/A _12997_/B vssd1 vssd1 vccd1 vccd1 _12998_/A sky130_fd_sc_hd__and2_1
XTAP_3671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_205_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17524_ _17544_/A _17524_/B vssd1 vssd1 vccd1 vccd1 _17524_/Y sky130_fd_sc_hd__nand2_1
XTAP_3693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14736_ _18310_/Q _18274_/Q _14736_/S vssd1 vssd1 vccd1 vccd1 _14736_/X sky130_fd_sc_hd__mux2_1
XFILLER_17_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11948_ _11980_/B vssd1 vssd1 vccd1 vccd1 _11948_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_1326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17455_ _18962_/Q _18926_/Q _17467_/S vssd1 vssd1 vccd1 vccd1 _17455_/X sky130_fd_sc_hd__mux2_1
XTAP_2992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14667_ _14681_/A _14670_/B vssd1 vssd1 vccd1 vccd1 _14667_/Y sky130_fd_sc_hd__nand2_1
X_11879_ _11879_/A _11879_/B vssd1 vssd1 vccd1 vccd1 _17832_/D sky130_fd_sc_hd__nor2_1
XFILLER_32_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16406_ _16524_/A vssd1 vssd1 vccd1 vccd1 _16450_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_177_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13618_ _14016_/A vssd1 vssd1 vccd1 vccd1 _13619_/A sky130_fd_sc_hd__buf_8
X_17386_ _18945_/Q _18909_/Q _17386_/S vssd1 vssd1 vccd1 vccd1 _17386_/X sky130_fd_sc_hd__mux2_1
XFILLER_158_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14598_ _14598_/A vssd1 vssd1 vccd1 vccd1 _14687_/A sky130_fd_sc_hd__buf_2
XFILLER_203_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_186_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_201_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16337_ _16521_/A vssd1 vssd1 vccd1 vccd1 _16389_/A sky130_fd_sc_hd__clkbuf_2
X_13549_ _13657_/A vssd1 vssd1 vccd1 vccd1 _13940_/A sky130_fd_sc_hd__buf_4
XFILLER_173_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_203_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_195_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_1280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16268_ _16268_/A _16268_/B vssd1 vssd1 vccd1 vccd1 _16268_/Y sky130_fd_sc_hd__nand2_1
XFILLER_145_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18007_ _18088_/CLK _18007_/D vssd1 vssd1 vccd1 vccd1 _18007_/Q sky130_fd_sc_hd__dfxtp_1
X_15219_ _18429_/Q _18393_/Q _15226_/S vssd1 vssd1 vccd1 vccd1 _15219_/X sky130_fd_sc_hd__mux2_1
X_16199_ _16199_/A _16202_/B vssd1 vssd1 vccd1 vccd1 _16199_/Y sky130_fd_sc_hd__nand2_1
XFILLER_12_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09711_ _09711_/A _09711_/B vssd1 vssd1 vccd1 vccd1 _09711_/X sky130_fd_sc_hd__or2_1
X_18909_ _18927_/CLK _18909_/D vssd1 vssd1 vccd1 vccd1 _18909_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_206_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09642_ _09664_/A _09642_/B vssd1 vssd1 vccd1 vccd1 _09649_/A sky130_fd_sc_hd__xor2_1
XFILLER_228_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19090__61 vssd1 vssd1 vccd1 vccd1 _19090__61/HI _19198_/A sky130_fd_sc_hd__conb_1
XFILLER_215_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09573_ _09573_/A _09573_/B vssd1 vssd1 vccd1 vccd1 _09573_/X sky130_fd_sc_hd__and2_1
XFILLER_222_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_230_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_223_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_208_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_211_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_221_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_221_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09007_ _09010_/A vssd1 vssd1 vccd1 vccd1 _09007_/Y sky130_fd_sc_hd__inv_2
XFILLER_151_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_219_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09909_ _10375_/S vssd1 vssd1 vccd1 vccd1 _09909_/X sky130_fd_sc_hd__buf_4
XFILLER_154_1290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12920_ _12920_/A _12920_/B _12920_/C vssd1 vssd1 vccd1 vccd1 _12921_/C sky130_fd_sc_hd__and3_1
XFILLER_4_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_207_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_207_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12851_ _17948_/Q _12851_/B vssd1 vssd1 vccd1 vccd1 _12852_/B sky130_fd_sc_hd__or2_1
XTAP_2211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11802_ _11930_/B vssd1 vssd1 vccd1 vccd1 _11976_/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15570_ _15570_/A _15570_/B vssd1 vssd1 vccd1 vccd1 _15570_/Y sky130_fd_sc_hd__nand2_1
XTAP_1510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12782_ _13019_/B _13041_/A vssd1 vssd1 vccd1 vccd1 _12783_/A sky130_fd_sc_hd__nand2_2
XTAP_2266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14521_ _18174_/Q _18173_/Q _18170_/Q _18169_/Q vssd1 vssd1 vccd1 vccd1 _14620_/A
+ sky130_fd_sc_hd__or4_2
XPHY_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11733_ _11742_/C vssd1 vssd1 vccd1 vccd1 _11733_/Y sky130_fd_sc_hd__inv_2
XTAP_1554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17240_ _17275_/A _17240_/B vssd1 vssd1 vccd1 vccd1 _17240_/Y sky130_fd_sc_hd__nand2_1
XFILLER_14_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14452_ _14452_/A _14452_/B vssd1 vssd1 vccd1 vccd1 _18203_/D sky130_fd_sc_hd__nor2_1
X_11664_ _11640_/Y _11651_/Y _11663_/X vssd1 vssd1 vccd1 vccd1 _11664_/X sky130_fd_sc_hd__a21o_1
XFILLER_109_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_202_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13403_ _10159_/A _11042_/X _11044_/B _11026_/A _13395_/X vssd1 vssd1 vccd1 vccd1
+ _18127_/D sky130_fd_sc_hd__o221a_1
XFILLER_211_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10615_ _10710_/B vssd1 vssd1 vccd1 vccd1 _12099_/A sky130_fd_sc_hd__clkbuf_4
X_17171_ _17458_/A _17202_/B vssd1 vssd1 vccd1 vccd1 _17180_/B sky130_fd_sc_hd__nor2_1
XFILLER_128_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14383_ _14383_/A _14383_/B _14383_/C vssd1 vssd1 vccd1 vccd1 _14384_/A sky130_fd_sc_hd__or3_1
X_11595_ _11595_/A _11681_/C vssd1 vssd1 vccd1 vccd1 _11595_/Y sky130_fd_sc_hd__nand2_1
XFILLER_183_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16122_ _18641_/Q _18605_/Q _16145_/S vssd1 vssd1 vccd1 vccd1 _16122_/X sky130_fd_sc_hd__mux2_1
XFILLER_167_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13334_ _14533_/A vssd1 vssd1 vccd1 vccd1 _13334_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_128_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10546_ _10536_/X _10538_/X _10541_/X _10545_/X _10939_/B _10903_/S vssd1 vssd1 vccd1
+ vccd1 _10547_/D sky130_fd_sc_hd__mux4_1
XFILLER_122_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16053_ _17265_/A _16366_/B vssd1 vssd1 vccd1 vccd1 _16127_/A sky130_fd_sc_hd__or2_1
XFILLER_183_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13265_ _13265_/A vssd1 vssd1 vccd1 vccd1 _18085_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_157_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10477_ _10935_/S _10477_/B vssd1 vssd1 vccd1 vccd1 _10477_/X sky130_fd_sc_hd__or2_1
X_15004_ _15083_/A vssd1 vssd1 vccd1 vccd1 _15004_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_12216_ _12216_/A vssd1 vssd1 vccd1 vccd1 _17853_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_29_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13196_ _13196_/A vssd1 vssd1 vccd1 vccd1 _18054_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_124_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12147_ _14457_/B vssd1 vssd1 vccd1 vccd1 _12147_/X sky130_fd_sc_hd__buf_6
XFILLER_150_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16955_ _16957_/B _16953_/X _16954_/Y _16940_/X vssd1 vssd1 vccd1 vccd1 _18802_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_133_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12078_ _12078_/A _12078_/B vssd1 vssd1 vccd1 vccd1 _12082_/A sky130_fd_sc_hd__xnor2_1
XFILLER_77_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15906_ _16055_/A _16043_/C vssd1 vssd1 vccd1 vccd1 _15913_/B sky130_fd_sc_hd__nor2_2
X_11029_ _17971_/Q _17970_/Q vssd1 vssd1 vccd1 vccd1 _11036_/B sky130_fd_sc_hd__and2_2
XFILLER_110_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16886_ _16886_/A vssd1 vssd1 vccd1 vccd1 _17480_/A sky130_fd_sc_hd__buf_4
XFILLER_77_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15837_ _15839_/B _15835_/X _15836_/Y _15823_/X vssd1 vssd1 vccd1 vccd1 _18538_/D
+ sky130_fd_sc_hd__o211a_1
X_18625_ _18658_/CLK _18625_/D vssd1 vssd1 vccd1 vccd1 _18625_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15768_ _15889_/A vssd1 vssd1 vccd1 vccd1 _15818_/A sky130_fd_sc_hd__clkbuf_2
X_18556_ _18557_/CLK _18556_/D vssd1 vssd1 vccd1 vccd1 _18556_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_212_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14719_ _18150_/Q _15015_/B vssd1 vssd1 vccd1 vccd1 _14833_/A sky130_fd_sc_hd__nand2_4
X_17507_ _17512_/B _17504_/X _17506_/X _17497_/X vssd1 vssd1 vccd1 vccd1 _18939_/D
+ sky130_fd_sc_hd__o211a_1
X_18487_ _18497_/CLK _18487_/D vssd1 vssd1 vccd1 vccd1 _18487_/Q sky130_fd_sc_hd__dfxtp_2
X_15699_ _15734_/A _15997_/B _15724_/C vssd1 vssd1 vccd1 vccd1 _15699_/X sky130_fd_sc_hd__or3_1
XFILLER_177_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17438_ _17444_/B _17436_/X _17437_/X _17421_/X vssd1 vssd1 vccd1 vccd1 _18921_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_178_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_220_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17369_ _17372_/B _17367_/X _17368_/Y _17361_/X vssd1 vssd1 vccd1 vccd1 _18904_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_146_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_68_wb_clk_i clkbuf_5_20_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18693_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_60_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_214_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_1346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09625_ _17974_/Q vssd1 vssd1 vccd1 vccd1 _10629_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_71_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09556_ _09560_/A _09591_/B vssd1 vssd1 vccd1 vccd1 _10038_/B sky130_fd_sc_hd__xnor2_4
XFILLER_231_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_1204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_197_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09487_ _13094_/A vssd1 vssd1 vccd1 vccd1 _12972_/A sky130_fd_sc_hd__buf_4
XFILLER_52_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_184_1283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_200_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_221_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_211_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_221_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10400_ _09349_/A _09354_/A _09344_/A _09349_/B _10349_/S _09937_/X vssd1 vssd1 vccd1
+ vccd1 _10400_/X sky130_fd_sc_hd__mux4_2
XFILLER_183_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11380_ _11368_/B _11297_/Y _11340_/B vssd1 vssd1 vccd1 vccd1 _11828_/B sky130_fd_sc_hd__o21ai_4
XFILLER_221_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_165_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10331_ _09237_/A _09227_/B _09232_/C _09237_/C _09958_/A _09948_/A vssd1 vssd1 vccd1
+ vccd1 _10331_/X sky130_fd_sc_hd__mux4_1
XFILLER_180_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13050_ _13050_/A vssd1 vssd1 vccd1 vccd1 _17995_/D sky130_fd_sc_hd__clkbuf_1
X_10262_ _10262_/A vssd1 vssd1 vccd1 vccd1 _10264_/A sky130_fd_sc_hd__clkinv_2
XFILLER_180_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12001_ _13438_/A _13426_/A vssd1 vssd1 vccd1 vccd1 _12026_/C sky130_fd_sc_hd__nand2_2
XFILLER_121_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10193_ _18120_/Q _10193_/B vssd1 vssd1 vccd1 vccd1 _10197_/A sky130_fd_sc_hd__xnor2_1
XFILLER_132_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19046__17 vssd1 vssd1 vccd1 vccd1 _19046__17/HI _19140_/A sky130_fd_sc_hd__conb_1
XFILLER_117_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_219_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16740_ _16760_/A vssd1 vssd1 vccd1 vccd1 _16740_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_59_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13952_ _18514_/Q _13738_/X _13950_/X _13951_/X vssd1 vssd1 vccd1 vccd1 _13952_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_4_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12903_ _17964_/Q _12904_/C _12902_/Y vssd1 vssd1 vccd1 vccd1 _17964_/D sky130_fd_sc_hd__a21oi_1
X_16671_ _18737_/Q _16670_/B _16670_/Y _16659_/X vssd1 vssd1 vccd1 vccd1 _18737_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_35_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13883_ _18880_/Q _13539_/A _13876_/X _13882_/X vssd1 vssd1 vccd1 vccd1 _13883_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_207_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18410_ _18443_/CLK _18410_/D vssd1 vssd1 vccd1 vccd1 _18410_/Q sky130_fd_sc_hd__dfxtp_2
X_15622_ _15736_/A vssd1 vssd1 vccd1 vccd1 _15717_/A sky130_fd_sc_hd__buf_2
XFILLER_46_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_185_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12834_ _12627_/B _12802_/Y _12832_/Y _17936_/Q _12833_/X vssd1 vssd1 vccd1 vccd1
+ _12835_/D sky130_fd_sc_hd__a221o_1
XTAP_2030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18341_ _18343_/CLK _18341_/D vssd1 vssd1 vccd1 vccd1 _18341_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15553_ _18505_/Q _18469_/Q _15565_/S vssd1 vssd1 vccd1 vccd1 _15553_/X sky130_fd_sc_hd__mux2_1
XFILLER_188_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12765_ _14373_/A _12762_/X _12764_/X vssd1 vssd1 vccd1 vccd1 _12765_/Y sky130_fd_sc_hd__o21ai_1
XTAP_2085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14504_ _18226_/Q _14504_/B vssd1 vssd1 vccd1 vccd1 _14505_/A sky130_fd_sc_hd__and2_1
XTAP_1373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18272_ _18275_/CLK _18272_/D vssd1 vssd1 vccd1 vccd1 _18272_/Q sky130_fd_sc_hd__dfxtp_1
X_11716_ _11716_/A _11716_/B vssd1 vssd1 vccd1 vccd1 _11860_/A sky130_fd_sc_hd__nand2_4
XTAP_1384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15484_ _15508_/A _15487_/B vssd1 vssd1 vccd1 vccd1 _15484_/Y sky130_fd_sc_hd__nand2_1
XTAP_1395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12696_ _17939_/Q _12697_/B vssd1 vssd1 vccd1 vccd1 _12698_/A sky130_fd_sc_hd__and2_1
XFILLER_30_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_175_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17223_ _17464_/A vssd1 vssd1 vccd1 vccd1 _17273_/A sky130_fd_sc_hd__clkbuf_2
X_14435_ _09501_/B _14405_/X _18199_/Q vssd1 vssd1 vccd1 vccd1 _14435_/X sky130_fd_sc_hd__o21a_1
X_11647_ _12251_/A _17861_/Q _11671_/B vssd1 vssd1 vccd1 vccd1 _12253_/A sky130_fd_sc_hd__nand3_2
XFILLER_156_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17154_ _17226_/A vssd1 vssd1 vccd1 vccd1 _17172_/S sky130_fd_sc_hd__buf_2
XFILLER_11_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14366_ _14381_/A vssd1 vssd1 vccd1 vccd1 _14366_/Y sky130_fd_sc_hd__inv_2
X_11578_ _11578_/A _11842_/A vssd1 vssd1 vccd1 vccd1 _11578_/Y sky130_fd_sc_hd__nand2_1
XFILLER_10_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16105_ _18637_/Q _18601_/Q _16113_/S vssd1 vssd1 vccd1 vccd1 _16105_/X sky130_fd_sc_hd__mux2_1
XFILLER_171_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13317_ _18091_/Q _18090_/Q vssd1 vssd1 vccd1 vccd1 _13317_/Y sky130_fd_sc_hd__nand2_1
X_10529_ _09165_/C _09170_/B _09160_/A _09160_/B _10484_/A _10489_/S vssd1 vssd1 vccd1
+ vccd1 _10529_/X sky130_fd_sc_hd__mux4_1
X_17085_ _17136_/A _17516_/B _17085_/C vssd1 vssd1 vccd1 vccd1 _17085_/X sky130_fd_sc_hd__or3_1
X_14297_ _14297_/A vssd1 vssd1 vccd1 vccd1 _14349_/A sky130_fd_sc_hd__buf_2
X_16036_ _16062_/A _16039_/B vssd1 vssd1 vccd1 vccd1 _16036_/Y sky130_fd_sc_hd__nand2_1
XFILLER_143_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13248_ _13248_/A vssd1 vssd1 vccd1 vccd1 _18077_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_83_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13179_ _13179_/A vssd1 vssd1 vccd1 vccd1 _18046_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_112_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17987_ _17987_/CLK _17987_/D vssd1 vssd1 vccd1 vccd1 _17987_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_112_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_211_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16938_ _18835_/Q _18799_/Q _16947_/S vssd1 vssd1 vccd1 vccd1 _16938_/X sky130_fd_sc_hd__mux2_1
XFILLER_226_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16869_ _18820_/Q _18784_/Q _16900_/S vssd1 vssd1 vccd1 vccd1 _16869_/X sky130_fd_sc_hd__mux2_1
XFILLER_20_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09410_ _18305_/Q _18304_/Q _18303_/Q vssd1 vssd1 vccd1 vccd1 _10956_/A sky130_fd_sc_hd__or3_4
XFILLER_16_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19060__31 vssd1 vssd1 vccd1 vccd1 _19060__31/HI _19154_/A sky130_fd_sc_hd__conb_1
X_18608_ _18608_/CLK _18608_/D vssd1 vssd1 vccd1 vccd1 _18608_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_129_1207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09341_ _18425_/Q _18424_/Q _18423_/Q vssd1 vssd1 vccd1 vccd1 _09344_/B sky130_fd_sc_hd__or3_4
X_18539_ _18542_/CLK _18539_/D vssd1 vssd1 vccd1 vccd1 _18539_/Q sky130_fd_sc_hd__dfxtp_2
Xclkbuf_leaf_186_wb_clk_i clkbuf_5_8_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17883_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_179_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09272_ _09272_/A _09440_/A vssd1 vssd1 vccd1 vccd1 _09435_/A sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_115_wb_clk_i clkbuf_5_31_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18467_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_221_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_166_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_159_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_1295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_138_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08987_ _08991_/A vssd1 vssd1 vccd1 vccd1 _08987_/Y sky130_fd_sc_hd__inv_2
XTAP_4905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_229_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_228_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09608_ _17982_/Q _09608_/B vssd1 vssd1 vccd1 vccd1 _09609_/B sky130_fd_sc_hd__xnor2_4
XFILLER_95_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10880_ _10757_/A _10875_/X _10879_/X _10833_/B vssd1 vssd1 vccd1 vccd1 _10880_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_3_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_231_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09539_ _18114_/Q vssd1 vssd1 vccd1 vccd1 _10181_/A sky130_fd_sc_hd__clkbuf_4
XPHY_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_189_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12550_ _17922_/Q vssd1 vssd1 vccd1 vccd1 _12564_/A sky130_fd_sc_hd__inv_2
XPHY_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11501_ _11501_/A _11501_/B _11501_/C _11500_/X vssd1 vssd1 vccd1 vccd1 _11501_/X
+ sky130_fd_sc_hd__or4b_4
XFILLER_106_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_200_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_197_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12481_ _17908_/Q _12499_/C vssd1 vssd1 vccd1 vccd1 _12484_/B sky130_fd_sc_hd__xor2_1
XFILLER_12_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14220_ _14349_/B _14342_/B vssd1 vssd1 vccd1 vccd1 _14323_/B sky130_fd_sc_hd__or2_1
X_11432_ _11419_/X _11431_/Y _11428_/B vssd1 vssd1 vccd1 vccd1 _11432_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_7_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14151_ _12019_/A _14135_/X _14142_/X _12019_/B _14150_/X vssd1 vssd1 vccd1 vccd1
+ _14151_/X sky130_fd_sc_hd__a221o_4
XFILLER_152_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11363_ _11404_/A _11307_/B _11403_/A vssd1 vssd1 vccd1 vccd1 _11364_/B sky130_fd_sc_hd__a21oi_1
X_13102_ _13102_/A vssd1 vssd1 vccd1 vccd1 _18011_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_3_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10314_ _09981_/X _10289_/Y _10312_/X _10313_/Y vssd1 vssd1 vccd1 vccd1 _10314_/X
+ sky130_fd_sc_hd__o211a_1
X_14082_ _18479_/Q _13617_/X _13619_/X _18455_/Q _14081_/X vssd1 vssd1 vccd1 vccd1
+ _14082_/X sky130_fd_sc_hd__a221o_1
X_11294_ _11951_/B vssd1 vssd1 vccd1 vccd1 _12023_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_98_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17910_ _17911_/CLK _17910_/D vssd1 vssd1 vccd1 vccd1 _17910_/Q sky130_fd_sc_hd__dfxtp_1
X_13033_ _13000_/B _13025_/X _13032_/X _13011_/X vssd1 vssd1 vccd1 vccd1 _17989_/D
+ sky130_fd_sc_hd__o211a_1
X_10245_ _09370_/C _09360_/D _09365_/B _09365_/D _10498_/A _12032_/A vssd1 vssd1 vccd1
+ vccd1 _10245_/X sky130_fd_sc_hd__mux4_2
XFILLER_79_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18890_ _18893_/CLK _18890_/D vssd1 vssd1 vccd1 vccd1 _18890_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_26_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17841_ _18157_/CLK _17841_/D vssd1 vssd1 vccd1 vccd1 _17841_/Q sky130_fd_sc_hd__dfxtp_1
X_10176_ _10422_/A vssd1 vssd1 vccd1 vccd1 _10939_/B sky130_fd_sc_hd__inv_2
XFILLER_67_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_226_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14984_ _14983_/B _14982_/X _14983_/Y _14980_/X vssd1 vssd1 vccd1 vccd1 _18335_/D
+ sky130_fd_sc_hd__o211a_1
X_17772_ _19030_/Q _12304_/Y _14436_/X vssd1 vssd1 vccd1 vccd1 _19030_/D sky130_fd_sc_hd__o21a_1
XFILLER_93_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_219_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16723_ _16755_/A _16723_/B vssd1 vssd1 vccd1 vccd1 _16723_/Y sky130_fd_sc_hd__nand2_1
X_13935_ _18325_/Q _13585_/A _13739_/X _18316_/Q vssd1 vssd1 vccd1 vccd1 _13935_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_207_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_228_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16654_ _18769_/Q _18733_/Q _16657_/S vssd1 vssd1 vccd1 vccd1 _16654_/X sky130_fd_sc_hd__mux2_1
X_13866_ _18841_/Q _13575_/X _13576_/X _18832_/Q _13865_/X vssd1 vssd1 vccd1 vccd1
+ _13866_/X sky130_fd_sc_hd__a221o_1
XFILLER_207_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15605_ _15633_/A _15605_/B vssd1 vssd1 vccd1 vccd1 _15605_/Y sky130_fd_sc_hd__nand2_1
XFILLER_90_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12817_ _12653_/B _17959_/Q _12796_/Y _17935_/Q vssd1 vssd1 vccd1 vccd1 _12817_/Y
+ sky130_fd_sc_hd__o22ai_1
X_16585_ _16631_/A _16589_/B vssd1 vssd1 vccd1 vccd1 _16585_/Y sky130_fd_sc_hd__nand2_1
XFILLER_22_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13797_ _18300_/Q _13759_/X _13780_/X _18291_/Q _13796_/X vssd1 vssd1 vccd1 vccd1
+ _13797_/X sky130_fd_sc_hd__a221o_4
XFILLER_15_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15536_ _15616_/A vssd1 vssd1 vccd1 vccd1 _15536_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_188_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18324_ _18324_/CLK _18324_/D vssd1 vssd1 vccd1 vccd1 _18324_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_37_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12748_ _12748_/A _12748_/B vssd1 vssd1 vccd1 vccd1 _12947_/A sky130_fd_sc_hd__or2_1
XFILLER_128_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_231_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_187_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18255_ _18266_/CLK _18255_/D vssd1 vssd1 vccd1 vccd1 _18255_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_147_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15467_ _15529_/A vssd1 vssd1 vccd1 vccd1 _15597_/B sky130_fd_sc_hd__buf_2
XFILLER_198_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12679_ _12679_/A _12679_/B vssd1 vssd1 vccd1 vccd1 _12679_/Y sky130_fd_sc_hd__nand2_1
XFILLER_8_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17206_ _17448_/A vssd1 vssd1 vccd1 vccd1 _17256_/A sky130_fd_sc_hd__buf_2
XFILLER_200_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14418_ _14404_/X _09497_/B _14405_/X vssd1 vssd1 vccd1 vccd1 _14418_/X sky130_fd_sc_hd__a21o_1
XFILLER_175_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18186_ _18230_/CLK _18186_/D vssd1 vssd1 vccd1 vccd1 _18186_/Q sky130_fd_sc_hd__dfxtp_1
X_15398_ _15403_/B _15395_/X _15397_/X _15382_/X vssd1 vssd1 vccd1 vccd1 _18432_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_191_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17137_ _17143_/B _17135_/X _17136_/X _17117_/X vssd1 vssd1 vccd1 vccd1 _18846_/D
+ sky130_fd_sc_hd__o211a_1
X_14349_ _14349_/A _14349_/B vssd1 vssd1 vccd1 vccd1 _14349_/Y sky130_fd_sc_hd__nand2_1
XFILLER_128_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17068_ _17091_/A _17068_/B vssd1 vssd1 vccd1 vccd1 _17068_/Y sky130_fd_sc_hd__nand2_1
XFILLER_170_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16019_ _16019_/A _16041_/B vssd1 vssd1 vccd1 vccd1 _16027_/B sky130_fd_sc_hd__nor2_2
XTAP_910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09890_ _18101_/Q _09918_/B vssd1 vssd1 vccd1 vccd1 _09915_/A sky130_fd_sc_hd__xnor2_4
XTAP_921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_214_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_211_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_214_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_226_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_230_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_213_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_230_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09324_ _18545_/Q _18544_/Q _18543_/Q vssd1 vssd1 vccd1 vccd1 _09327_/B sky130_fd_sc_hd__or3_2
XFILLER_55_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_222_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_178_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09255_ _09255_/A _09254_/Y vssd1 vssd1 vccd1 vccd1 _09272_/A sky130_fd_sc_hd__or2b_1
XFILLER_107_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_222_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09186_ _09186_/A _09186_/B _09186_/C _09186_/D vssd1 vssd1 vccd1 vccd1 _09187_/C
+ sky130_fd_sc_hd__and4_1
XFILLER_88_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_181_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_83_wb_clk_i clkbuf_5_23_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18614_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_161_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_12_wb_clk_i clkbuf_5_4_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17965_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_89_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10030_ _09720_/A _10022_/X _10029_/X _09657_/A vssd1 vssd1 vccd1 vccd1 _10030_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_5414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11981_ _11968_/X _11978_/X _12022_/B vssd1 vssd1 vccd1 vccd1 _13421_/A sky130_fd_sc_hd__a21oi_2
XFILLER_75_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13720_ _13720_/A vssd1 vssd1 vccd1 vccd1 _13721_/A sky130_fd_sc_hd__buf_6
XFILLER_29_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10932_ _10932_/A _10932_/B vssd1 vssd1 vccd1 vccd1 _10932_/X sky130_fd_sc_hd__and2_1
XFILLER_216_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_204_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_216_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13651_ _13733_/A vssd1 vssd1 vccd1 vccd1 _13651_/X sky130_fd_sc_hd__buf_6
X_10863_ _10910_/C _10861_/X _10862_/X _10843_/X vssd1 vssd1 vccd1 vccd1 _10863_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_220_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_213_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12602_ _12597_/B _12529_/X _11218_/X vssd1 vssd1 vccd1 vccd1 _12602_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_71_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16370_ _16501_/B vssd1 vssd1 vccd1 vccd1 _16422_/C sky130_fd_sc_hd__clkbuf_2
XPHY_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13582_ _13582_/A vssd1 vssd1 vccd1 vccd1 _13582_/X sky130_fd_sc_hd__buf_6
XFILLER_73_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10794_ _09219_/A _09209_/C _10812_/S vssd1 vssd1 vccd1 vccd1 _10794_/X sky130_fd_sc_hd__mux2_1
XPHY_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15321_ _15325_/B _15317_/X _15320_/Y _15315_/X vssd1 vssd1 vccd1 vccd1 _18415_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_158_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12533_ _17917_/Q vssd1 vssd1 vccd1 vccd1 _12533_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_160_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_201_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18040_ _18094_/CLK _18040_/D vssd1 vssd1 vccd1 vccd1 _18040_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_40_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15252_ _15252_/A vssd1 vssd1 vccd1 vccd1 _15303_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_12_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12464_ _17905_/Q _12470_/B vssd1 vssd1 vccd1 vccd1 _12477_/C sky130_fd_sc_hd__xor2_2
XFILLER_200_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_201_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14203_ _14297_/A vssd1 vssd1 vccd1 vccd1 _14203_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_125_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11415_ _19029_/Q _11415_/B vssd1 vssd1 vccd1 vccd1 _11415_/Y sky130_fd_sc_hd__nand2_1
XFILLER_32_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15183_ _15182_/B _15181_/X _15182_/Y _15166_/X vssd1 vssd1 vccd1 vccd1 _18383_/D
+ sky130_fd_sc_hd__o211a_1
X_12395_ _12406_/A _12395_/B vssd1 vssd1 vccd1 vccd1 _12397_/C sky130_fd_sc_hd__nor2_1
XFILLER_158_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_153_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14134_ _18275_/Q _13546_/A _14130_/X _14133_/X vssd1 vssd1 vccd1 vccd1 _14134_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_126_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11346_ _11346_/A _11388_/A vssd1 vssd1 vccd1 vccd1 _11346_/Y sky130_fd_sc_hd__nand2_1
XFILLER_4_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_152_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14065_ _12028_/A _14057_/X _14064_/X _12055_/B vssd1 vssd1 vccd1 vccd1 _14065_/X
+ sky130_fd_sc_hd__a22o_1
X_18942_ _18953_/CLK _18942_/D vssd1 vssd1 vccd1 vccd1 _18942_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_165_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11277_ _11281_/A _12041_/A _11277_/C vssd1 vssd1 vccd1 vccd1 _11812_/B sky130_fd_sc_hd__or3_1
X_13016_ _18151_/Q vssd1 vssd1 vccd1 vccd1 _13016_/X sky130_fd_sc_hd__buf_2
X_10228_ _10560_/S vssd1 vssd1 vccd1 vccd1 _10559_/S sky130_fd_sc_hd__clkbuf_2
X_18873_ _18875_/CLK _18873_/D vssd1 vssd1 vccd1 vccd1 _18873_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_121_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_228_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17824_ _17824_/CLK _17824_/D vssd1 vssd1 vccd1 vccd1 _17824_/Q sky130_fd_sc_hd__dfxtp_1
Xhold2 hold2/A vssd1 vssd1 vccd1 vccd1 hold2/X sky130_fd_sc_hd__clkdlybuf4s50_1
X_10159_ _10159_/A _10159_/B vssd1 vssd1 vccd1 vccd1 _10162_/A sky130_fd_sc_hd__xnor2_1
XFILLER_67_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_227_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_181_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14967_ _18367_/Q _18331_/Q _14974_/S vssd1 vssd1 vccd1 vccd1 _14967_/X sky130_fd_sc_hd__mux2_1
X_17755_ _17755_/A vssd1 vssd1 vccd1 vccd1 _19020_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_54_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16706_ _18781_/Q _18745_/Q _16715_/S vssd1 vssd1 vccd1 vccd1 _16706_/X sky130_fd_sc_hd__mux2_1
XFILLER_78_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13918_ _18757_/Q _13856_/A _13588_/X _18748_/Q _13917_/X vssd1 vssd1 vccd1 vccd1
+ _13918_/X sky130_fd_sc_hd__a221o_1
XFILLER_130_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14898_ _14900_/B _14896_/X _14897_/Y _14881_/X vssd1 vssd1 vccd1 vccd1 _18313_/D
+ sky130_fd_sc_hd__o211a_1
X_17686_ _17686_/A vssd1 vssd1 vccd1 vccd1 _18983_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_208_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_1278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13849_ _18721_/Q _13848_/X _13588_/X _18712_/Q vssd1 vssd1 vccd1 vccd1 _13849_/X
+ sky130_fd_sc_hd__a22o_1
X_16637_ _18765_/Q _18729_/Q _16637_/S vssd1 vssd1 vccd1 vccd1 _16637_/X sky130_fd_sc_hd__mux2_1
XFILLER_23_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_223_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16568_ _16615_/A _16716_/B _16568_/C vssd1 vssd1 vccd1 vccd1 _16568_/X sky130_fd_sc_hd__or3_1
XFILLER_222_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_210_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18307_ _18307_/CLK _18307_/D vssd1 vssd1 vccd1 vccd1 _18307_/Q sky130_fd_sc_hd__dfxtp_2
X_15519_ _18496_/Q _18460_/Q _15545_/S vssd1 vssd1 vccd1 vccd1 _15519_/X sky130_fd_sc_hd__mux2_1
XFILLER_200_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16499_ _16510_/A _16499_/B vssd1 vssd1 vccd1 vccd1 _16499_/Y sky130_fd_sc_hd__nand2_1
XFILLER_175_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09040_ _09040_/A vssd1 vssd1 vccd1 vccd1 _09040_/Y sky130_fd_sc_hd__inv_2
XFILLER_175_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18238_ _18263_/CLK _18238_/D vssd1 vssd1 vccd1 vccd1 _18238_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_191_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18169_ _18184_/CLK _18169_/D vssd1 vssd1 vccd1 vccd1 _18169_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_128_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_1366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09942_ _09974_/A vssd1 vssd1 vccd1 vccd1 _10333_/S sky130_fd_sc_hd__clkbuf_4
XTAP_740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09873_ _09876_/A _09876_/B _09872_/Y vssd1 vssd1 vccd1 vccd1 _09880_/A sky130_fd_sc_hd__o21ba_1
XTAP_751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_225_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_15 _09176_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_26 _09253_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_37 _12123_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XINSDIODE2_48 _10500_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_59 _14457_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_1338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_130_wb_clk_i clkbuf_5_25_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18404_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_53_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_213_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09307_ _18458_/Q _18457_/Q _18456_/Q vssd1 vssd1 vccd1 vccd1 _09309_/C sky130_fd_sc_hd__or3_2
XFILLER_70_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_210_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09238_ _09238_/A _09238_/B _09238_/C vssd1 vssd1 vccd1 vccd1 _09255_/A sky130_fd_sc_hd__and3_2
XFILLER_6_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09169_ _18635_/Q _18634_/Q _18633_/Q vssd1 vssd1 vccd1 vccd1 _09170_/D sky130_fd_sc_hd__or3_4
XFILLER_108_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11200_ _11201_/A _11205_/C vssd1 vssd1 vccd1 vccd1 _11202_/B sky130_fd_sc_hd__or2_1
XFILLER_108_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12180_ _12180_/A _12180_/B vssd1 vssd1 vccd1 vccd1 _12180_/Y sky130_fd_sc_hd__nor2_1
XFILLER_79_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_218_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11131_ _11541_/A vssd1 vssd1 vccd1 vccd1 _11453_/A sky130_fd_sc_hd__buf_2
XFILLER_218_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11062_ _17817_/Q vssd1 vssd1 vccd1 vccd1 _11224_/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_5211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_1216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10013_ _10060_/A vssd1 vssd1 vccd1 vccd1 _10096_/S sky130_fd_sc_hd__buf_4
XTAP_5244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15870_ _15921_/A _16021_/B _15870_/C vssd1 vssd1 vccd1 vccd1 _15870_/X sky130_fd_sc_hd__or3_1
XFILLER_95_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_218_wb_clk_i _17864_/CLK vssd1 vssd1 vccd1 vccd1 _19031_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_5266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14821_ _18331_/Q _18295_/Q _14830_/S vssd1 vssd1 vccd1 vccd1 _14821_/X sky130_fd_sc_hd__mux2_1
XFILLER_36_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_218_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_229_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14752_ _18314_/Q _18278_/Q _14756_/S vssd1 vssd1 vccd1 vccd1 _14752_/X sky130_fd_sc_hd__mux2_1
X_17540_ _18985_/Q _18949_/Q _17543_/S vssd1 vssd1 vccd1 vccd1 _17540_/X sky130_fd_sc_hd__mux2_1
XTAP_3864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11964_ _11964_/A _12015_/A _11964_/C _12026_/D vssd1 vssd1 vccd1 vccd1 _12020_/B
+ sky130_fd_sc_hd__and4_1
XTAP_3875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_229_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13703_ _13703_/A vssd1 vssd1 vccd1 vccd1 _14030_/A sky130_fd_sc_hd__buf_4
XTAP_3886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10915_ _09319_/D _09309_/D _09309_/A _10575_/A _10498_/A _12032_/A vssd1 vssd1 vccd1
+ vccd1 _10915_/X sky130_fd_sc_hd__mux4_1
XTAP_3897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17471_ _17471_/A _17538_/C vssd1 vssd1 vccd1 vccd1 _17477_/B sky130_fd_sc_hd__nor2_1
X_14683_ _14683_/A _14683_/B vssd1 vssd1 vccd1 vccd1 _14683_/Y sky130_fd_sc_hd__nand2_1
XFILLER_60_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11895_ _11895_/A vssd1 vssd1 vccd1 vccd1 _14457_/B sky130_fd_sc_hd__buf_6
XFILLER_229_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19210_ _19210_/A _08979_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[10] sky130_fd_sc_hd__ebufn_8
X_16422_ _16434_/A _16716_/B _16422_/C vssd1 vssd1 vccd1 vccd1 _16422_/X sky130_fd_sc_hd__or3_1
X_13634_ _18480_/Q _13612_/X _13620_/X _13633_/X vssd1 vssd1 vccd1 vccd1 _13634_/X
+ sky130_fd_sc_hd__a211o_2
X_10846_ _10829_/X _10845_/X _10757_/A vssd1 vssd1 vccd1 vccd1 _10846_/X sky130_fd_sc_hd__a21o_1
XFILLER_32_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_204_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_198_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16353_ _16392_/A _16353_/B vssd1 vssd1 vccd1 vccd1 _16353_/Y sky130_fd_sc_hd__nand2_1
X_19141_ _19141_/A _09055_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[11] sky130_fd_sc_hd__ebufn_8
X_13565_ _13715_/A vssd1 vssd1 vccd1 vccd1 _13566_/A sky130_fd_sc_hd__buf_6
XFILLER_160_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10777_ _10779_/A _10777_/B vssd1 vssd1 vccd1 vccd1 _10777_/X sky130_fd_sc_hd__or2_1
XFILLER_73_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_200_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15304_ _18413_/Q _15303_/B _15303_/Y _15283_/X vssd1 vssd1 vccd1 vccd1 _18413_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_157_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12516_ _11763_/A _11763_/C _12514_/Y _17543_/S _11767_/B vssd1 vssd1 vccd1 vccd1
+ _12517_/B sky130_fd_sc_hd__a32o_1
X_16284_ _16524_/A vssd1 vssd1 vccd1 vccd1 _16329_/A sky130_fd_sc_hd__buf_2
XFILLER_158_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13496_ _13720_/A vssd1 vssd1 vccd1 vccd1 _13763_/A sky130_fd_sc_hd__buf_6
XFILLER_125_1298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15235_ _18433_/Q _18397_/Q _15246_/S vssd1 vssd1 vccd1 vccd1 _15235_/X sky130_fd_sc_hd__mux2_1
X_18023_ _18030_/CLK _18023_/D vssd1 vssd1 vccd1 vccd1 _18023_/Q sky130_fd_sc_hd__dfxtp_1
X_12447_ _12452_/A _12444_/Y _12437_/A _12438_/Y vssd1 vssd1 vccd1 vccd1 _12447_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_172_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15166_ _15187_/A vssd1 vssd1 vccd1 vccd1 _15166_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_5_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12378_ _12388_/A _12375_/Y _12365_/X _12369_/B vssd1 vssd1 vccd1 vccd1 _12379_/C
+ sky130_fd_sc_hd__o211ai_1
XFILLER_181_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14117_ _18926_/Q _13515_/X _13500_/X _18944_/Q vssd1 vssd1 vccd1 vccd1 _14117_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_158_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11329_ _17877_/Q _11339_/C _11385_/B vssd1 vssd1 vccd1 vccd1 _11329_/Y sky130_fd_sc_hd__nand3_1
X_15097_ _18399_/Q _18363_/Q _15100_/S vssd1 vssd1 vccd1 vccd1 _15097_/X sky130_fd_sc_hd__mux2_1
XFILLER_119_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14048_ _18539_/Q _13524_/A _13621_/A _18542_/Q _14047_/X vssd1 vssd1 vccd1 vccd1
+ _14048_/X sky130_fd_sc_hd__a221o_1
XFILLER_141_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18925_ _18926_/CLK _18925_/D vssd1 vssd1 vccd1 vccd1 _18925_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_80_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18856_ _18862_/CLK _18856_/D vssd1 vssd1 vccd1 vccd1 _18856_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_68_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_227_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17807_ _18191_/CLK _17807_/D vssd1 vssd1 vccd1 vccd1 _17807_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_55_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18787_ _18788_/CLK _18787_/D vssd1 vssd1 vccd1 vccd1 _18787_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_55_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15999_ _18613_/Q _18577_/Q _16010_/S vssd1 vssd1 vccd1 vccd1 _15999_/X sky130_fd_sc_hd__mux2_1
X_17738_ _17738_/A vssd1 vssd1 vccd1 vccd1 _19012_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_224_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINSDIODE2_130 _16431_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17669_ _17681_/A _17669_/B vssd1 vssd1 vccd1 vccd1 _17670_/A sky130_fd_sc_hd__and2_1
XFILLER_208_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_141 _17265_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XINSDIODE2_152 _18420_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XINSDIODE2_163 _18360_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_174 _18705_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_211_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_185 _09098_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_1321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_196 _10795_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09023_ _09029_/A vssd1 vssd1 vccd1 vccd1 _09028_/A sky130_fd_sc_hd__buf_12
XFILLER_156_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09925_ _10376_/B vssd1 vssd1 vccd1 vccd1 _12124_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_59_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09856_ _09858_/B _09858_/A vssd1 vssd1 vccd1 vccd1 _09860_/B sky130_fd_sc_hd__and2b_1
XFILLER_112_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_219_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09787_ _09787_/A _09787_/B vssd1 vssd1 vccd1 vccd1 _09793_/B sky130_fd_sc_hd__xnor2_1
XTAP_3116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_215_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_198_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10700_ _10694_/X _10697_/X _10700_/S vssd1 vssd1 vccd1 vccd1 _10700_/X sky130_fd_sc_hd__mux2_1
XTAP_1747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11680_ _11680_/A _11850_/A _11680_/C _11680_/D vssd1 vssd1 vccd1 vccd1 _11716_/A
+ sky130_fd_sc_hd__or4_1
XFILLER_41_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_201_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10631_ _10661_/A _10661_/B _10630_/X vssd1 vssd1 vccd1 vccd1 _10650_/B sky130_fd_sc_hd__a21o_4
XFILLER_41_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_220_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_195_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13350_ _18101_/Q _13336_/X _11023_/X vssd1 vssd1 vccd1 vccd1 _18101_/D sky130_fd_sc_hd__o21a_1
XFILLER_224_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10562_ _09198_/C _09203_/D _09203_/A _09193_/D _10494_/A _10462_/X vssd1 vssd1 vccd1
+ vccd1 _10562_/X sky130_fd_sc_hd__mux4_1
XFILLER_14_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12301_ _12301_/A vssd1 vssd1 vccd1 vccd1 _12301_/Y sky130_fd_sc_hd__inv_2
X_13281_ _13281_/A _13281_/B vssd1 vssd1 vccd1 vccd1 _13292_/B sky130_fd_sc_hd__or2_1
X_10493_ _10419_/A _10488_/X _10492_/X _10270_/A vssd1 vssd1 vccd1 vccd1 _10493_/X
+ sky130_fd_sc_hd__o211a_1
X_15020_ _15025_/B _15018_/X _15019_/X _15004_/X vssd1 vssd1 vccd1 vccd1 _18342_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_136_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12232_ _11614_/A _12221_/A _12233_/A vssd1 vssd1 vccd1 vccd1 _12232_/X sky130_fd_sc_hd__a21o_1
XFILLER_120_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12163_ _14436_/A vssd1 vssd1 vccd1 vccd1 _12163_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_68_1277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_150_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11114_ _11114_/A vssd1 vssd1 vccd1 vccd1 _17797_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_155_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16971_ _17168_/A vssd1 vssd1 vccd1 vccd1 _17035_/A sky130_fd_sc_hd__buf_2
X_12094_ _12094_/A _13494_/B vssd1 vssd1 vccd1 vccd1 _12095_/D sky130_fd_sc_hd__xnor2_1
XFILLER_89_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18710_ _18710_/CLK _18710_/D vssd1 vssd1 vccd1 vccd1 _18710_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_1_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15922_ _15928_/B _15920_/X _15921_/X _15901_/X vssd1 vssd1 vccd1 vccd1 _18558_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_5030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11045_ _13346_/A vssd1 vssd1 vccd1 vccd1 _11045_/X sky130_fd_sc_hd__clkbuf_2
XTAP_5041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18641_ _18641_/CLK _18641_/D vssd1 vssd1 vccd1 vccd1 _18641_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_209_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15853_ _15876_/A _15853_/B vssd1 vssd1 vccd1 vccd1 _15853_/Y sky130_fd_sc_hd__nand2_1
XTAP_5085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14804_ _15241_/A _14841_/B vssd1 vssd1 vccd1 vccd1 _14814_/B sky130_fd_sc_hd__nor2_2
XFILLER_91_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18572_ _18572_/CLK _18572_/D vssd1 vssd1 vccd1 vccd1 _18572_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_4384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15784_ _15782_/B _15781_/X _15782_/Y _15783_/X vssd1 vssd1 vccd1 vccd1 _18524_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_4395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12996_ _12991_/X _12994_/X _12995_/X _13000_/B vssd1 vssd1 vccd1 vccd1 _12997_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_166_1310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17523_ _18980_/Q _18944_/Q _17533_/S vssd1 vssd1 vccd1 vccd1 _17523_/X sky130_fd_sc_hd__mux2_1
XFILLER_91_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_189_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14735_ _14742_/B _14733_/X _14734_/X _14716_/X vssd1 vssd1 vccd1 vccd1 _18273_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_45_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11947_ _11947_/A _11947_/B vssd1 vssd1 vccd1 vccd1 _11980_/B sky130_fd_sc_hd__and2_1
XTAP_3694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14666_ _18258_/Q _14670_/B _14665_/X _14647_/X vssd1 vssd1 vccd1 vccd1 _18258_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_60_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17454_ _17456_/B _17452_/X _17453_/Y _17441_/X vssd1 vssd1 vccd1 vccd1 _18925_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_2993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_1338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11878_ hold2/X _11867_/X _11875_/Y vssd1 vssd1 vccd1 vccd1 _11879_/B sky130_fd_sc_hd__a21oi_1
XFILLER_221_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16405_ _18707_/Q _18671_/Q _16421_/S vssd1 vssd1 vccd1 vccd1 _16405_/X sky130_fd_sc_hd__mux2_1
X_13617_ _13617_/A vssd1 vssd1 vccd1 vccd1 _13617_/X sky130_fd_sc_hd__buf_6
X_10829_ _10829_/A vssd1 vssd1 vccd1 vccd1 _10829_/X sky130_fd_sc_hd__buf_4
XFILLER_220_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14597_ _14597_/A vssd1 vssd1 vccd1 vccd1 _14665_/A sky130_fd_sc_hd__clkbuf_4
X_17385_ _17526_/A _17397_/B vssd1 vssd1 vccd1 vccd1 _17395_/B sky130_fd_sc_hd__nor2_1
XFILLER_119_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16336_ _18691_/Q _18655_/Q _16345_/S vssd1 vssd1 vccd1 vccd1 _16336_/X sky130_fd_sc_hd__mux2_1
X_13548_ _13613_/A vssd1 vssd1 vccd1 vccd1 _13657_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_119_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16267_ _18674_/Q _18638_/Q _16271_/S vssd1 vssd1 vccd1 vccd1 _16267_/X sky130_fd_sc_hd__mux2_1
XFILLER_145_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13479_ _17847_/Q _13457_/A _13465_/A vssd1 vssd1 vccd1 vccd1 _13480_/B sky130_fd_sc_hd__a21oi_1
XFILLER_199_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15218_ _15218_/A _15229_/B vssd1 vssd1 vccd1 vccd1 _15227_/B sky130_fd_sc_hd__nor2_2
XFILLER_161_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18006_ _18088_/CLK _18006_/D vssd1 vssd1 vccd1 vccd1 _18006_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_145_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16198_ _18658_/Q _18622_/Q _16215_/S vssd1 vssd1 vccd1 vccd1 _16198_/X sky130_fd_sc_hd__mux2_1
XFILLER_161_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15149_ _15277_/B vssd1 vssd1 vccd1 vccd1 _15199_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_113_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_214_1333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_206_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09710_ _09695_/X _09696_/X _09697_/X _09698_/X _10942_/A _09709_/X vssd1 vssd1 vccd1
+ vccd1 _09711_/B sky130_fd_sc_hd__mux4_1
X_18908_ _18908_/CLK _18908_/D vssd1 vssd1 vccd1 vccd1 _18908_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_132_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09641_ _09668_/A vssd1 vssd1 vccd1 vccd1 _12078_/A sky130_fd_sc_hd__buf_4
X_18839_ _18845_/CLK _18839_/D vssd1 vssd1 vccd1 vccd1 _18839_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_83_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_222_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09572_ _09573_/A _09573_/B vssd1 vssd1 vccd1 vccd1 _09592_/B sky130_fd_sc_hd__xor2_1
XFILLER_83_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_209_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_209_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_222_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_212_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_223_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_196_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_180_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_211_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_195_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_221_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_177_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09006_ _09010_/A vssd1 vssd1 vccd1 vccd1 _09006_/Y sky130_fd_sc_hd__inv_2
XFILLER_152_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_219_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_215_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09908_ _10348_/A vssd1 vssd1 vccd1 vccd1 _10375_/S sky130_fd_sc_hd__buf_2
XFILLER_219_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09839_ _09839_/A _09840_/B vssd1 vssd1 vccd1 vccd1 _09855_/B sky130_fd_sc_hd__xor2_4
XFILLER_111_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12850_ _17948_/Q _12851_/B vssd1 vssd1 vccd1 vccd1 _12857_/C sky130_fd_sc_hd__and2_1
XFILLER_74_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11801_ _17789_/Q _17788_/Q _17790_/Q vssd1 vssd1 vccd1 vccd1 _11930_/B sky130_fd_sc_hd__o21ai_2
XFILLER_215_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12781_ _18152_/Q _12781_/B vssd1 vssd1 vccd1 vccd1 _13041_/A sky130_fd_sc_hd__nor2_2
XTAP_2245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_3_1_0_wb_clk_i clkbuf_3_1_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_4_3_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_14_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14520_ _18172_/Q _18171_/Q vssd1 vssd1 vccd1 vccd1 _14593_/A sky130_fd_sc_hd__or2_1
XFILLER_202_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11732_ _11732_/A _11732_/B vssd1 vssd1 vccd1 vccd1 _11742_/C sky130_fd_sc_hd__xnor2_1
XTAP_1544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14451_ _18203_/Q _14450_/Y _14428_/X _09505_/B vssd1 vssd1 vccd1 vccd1 _14452_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_109_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11663_ _11683_/B _11663_/B _11683_/A vssd1 vssd1 vccd1 vccd1 _11663_/X sky130_fd_sc_hd__or3b_1
XTAP_1599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13402_ _13402_/A vssd1 vssd1 vccd1 vccd1 _18126_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_174_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10614_ _10731_/B _10614_/B vssd1 vssd1 vccd1 vccd1 _10710_/B sky130_fd_sc_hd__or2_1
X_17170_ _17169_/B _17167_/X _17169_/Y _17161_/X vssd1 vssd1 vccd1 vccd1 _18854_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_161_1262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14382_ _14379_/Y _14381_/X _17766_/A vssd1 vssd1 vccd1 vccd1 _18188_/D sky130_fd_sc_hd__a21oi_1
XFILLER_195_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11594_ _11594_/A vssd1 vssd1 vccd1 vccd1 _11681_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_35_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16121_ _16123_/B _16118_/X _16119_/Y _16120_/X vssd1 vssd1 vccd1 vccd1 _18604_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_195_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13333_ _13318_/A _13318_/B _13332_/Y _13324_/A vssd1 vssd1 vccd1 vccd1 _13333_/Y
+ sky130_fd_sc_hd__o31ai_1
XFILLER_70_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10545_ _10543_/X _10544_/X _10549_/A vssd1 vssd1 vccd1 vccd1 _10545_/X sky130_fd_sc_hd__mux2_1
XFILLER_183_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16052_ _16051_/B _16050_/X _16051_/Y _16048_/X vssd1 vssd1 vccd1 vccd1 _18590_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_170_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13264_ _13266_/A _18086_/Q vssd1 vssd1 vccd1 vccd1 _13265_/A sky130_fd_sc_hd__and2_1
XFILLER_196_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10476_ _09248_/B _09243_/B _09253_/C _09243_/C _10412_/A _10411_/A vssd1 vssd1 vccd1
+ vccd1 _10477_/B sky130_fd_sc_hd__mux4_1
XFILLER_182_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15003_ _15207_/A vssd1 vssd1 vccd1 vccd1 _15083_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_136_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12215_ _14504_/B _12239_/C _12215_/C vssd1 vssd1 vccd1 vccd1 _12216_/A sky130_fd_sc_hd__and3_1
XFILLER_108_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13195_ _13197_/A _18055_/Q vssd1 vssd1 vccd1 vccd1 _13196_/A sky130_fd_sc_hd__and2_1
XFILLER_29_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12146_ _12183_/B _12158_/A _12169_/B vssd1 vssd1 vccd1 vccd1 _12146_/X sky130_fd_sc_hd__or3_1
XFILLER_150_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16954_ _16954_/A _16957_/B vssd1 vssd1 vccd1 vccd1 _16954_/Y sky130_fd_sc_hd__nand2_1
XFILLER_81_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12077_ _17977_/Q _12077_/B vssd1 vssd1 vccd1 vccd1 _12078_/B sky130_fd_sc_hd__xnor2_1
XFILLER_38_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15905_ _15975_/A vssd1 vssd1 vccd1 vccd1 _16043_/C sky130_fd_sc_hd__buf_2
X_11028_ _17971_/Q _17970_/Q vssd1 vssd1 vccd1 vccd1 _11031_/A sky130_fd_sc_hd__nor2_1
XFILLER_37_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16885_ _18788_/Q _16884_/B _16884_/Y _16871_/X vssd1 vssd1 vccd1 vccd1 _18788_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_2_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_225_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18624_ _18658_/CLK _18624_/D vssd1 vssd1 vccd1 vccd1 _18624_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_49_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15836_ _15873_/A _15839_/B vssd1 vssd1 vccd1 vccd1 _15836_/Y sky130_fd_sc_hd__nand2_1
XTAP_4170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18555_ _18557_/CLK _18555_/D vssd1 vssd1 vccd1 vccd1 _18555_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_24_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15767_ _18520_/Q _15769_/B _15766_/Y _15763_/X vssd1 vssd1 vccd1 vccd1 _18520_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_3480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12979_ _12975_/A _12952_/X _12978_/X _12964_/X vssd1 vssd1 vccd1 vccd1 _17976_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_206_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17506_ _17538_/A _17506_/B _17516_/C vssd1 vssd1 vccd1 vccd1 _17506_/X sky130_fd_sc_hd__or3_1
XFILLER_206_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14718_ _15156_/A _14843_/C vssd1 vssd1 vccd1 vccd1 _14729_/B sky130_fd_sc_hd__nor2_2
XFILLER_127_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18486_ _18497_/CLK _18486_/D vssd1 vssd1 vccd1 vccd1 _18486_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_75_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15698_ _18540_/Q _18504_/Q _15714_/S vssd1 vssd1 vccd1 vccd1 _15698_/X sky130_fd_sc_hd__mux2_1
XTAP_2790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_220_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17437_ _17437_/A _17437_/B _17460_/C vssd1 vssd1 vccd1 vccd1 _17437_/X sky130_fd_sc_hd__or3_1
X_14649_ _17674_/A _14660_/B vssd1 vssd1 vccd1 vccd1 _16919_/A sky130_fd_sc_hd__or2_4
XFILLER_60_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_220_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_221_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_193_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17368_ _17392_/A _17372_/B vssd1 vssd1 vccd1 vccd1 _17368_/Y sky130_fd_sc_hd__nand2_1
XFILLER_159_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16319_ _16757_/A _16356_/B vssd1 vssd1 vccd1 vccd1 _16329_/B sky130_fd_sc_hd__nor2_2
XFILLER_192_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_173_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17299_ _17334_/A _17303_/B vssd1 vssd1 vccd1 vccd1 _17299_/Y sky130_fd_sc_hd__nand2_1
XFILLER_146_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_229_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_228_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_214_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_228_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09624_ _09645_/A vssd1 vssd1 vccd1 vccd1 _13372_/A sky130_fd_sc_hd__buf_2
XFILLER_3_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09555_ _09590_/B _09555_/B vssd1 vssd1 vccd1 vccd1 _09591_/B sky130_fd_sc_hd__xnor2_4
XFILLER_71_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_37_wb_clk_i clkbuf_5_18_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18806_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_43_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_212_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09486_ _12224_/A vssd1 vssd1 vccd1 vccd1 _13094_/A sky130_fd_sc_hd__buf_2
XFILLER_58_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_212_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_1295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_225_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_196_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_221_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_221_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10330_ _09227_/C _09232_/B _09237_/D _09232_/D _10285_/S _09959_/X vssd1 vssd1 vccd1
+ vccd1 _10330_/X sky130_fd_sc_hd__mux4_2
XFILLER_125_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_124_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10261_ _11910_/A _11910_/B vssd1 vssd1 vccd1 vccd1 _10262_/A sky130_fd_sc_hd__xnor2_1
XFILLER_191_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12000_ _12006_/A _12006_/B _11973_/B vssd1 vssd1 vccd1 vccd1 _12019_/A sky130_fd_sc_hd__a21oi_4
XFILLER_191_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10192_ _10215_/A _10192_/B vssd1 vssd1 vccd1 vccd1 _10246_/A sky130_fd_sc_hd__xnor2_1
XFILLER_121_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_219_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13951_ _18502_/Q _13742_/X _13743_/X _18484_/Q vssd1 vssd1 vccd1 vccd1 _13951_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_120_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12902_ _17964_/Q _12904_/C _12874_/X vssd1 vssd1 vccd1 vccd1 _12902_/Y sky130_fd_sc_hd__o21ai_1
X_16670_ _16699_/A _16670_/B vssd1 vssd1 vccd1 vccd1 _16670_/Y sky130_fd_sc_hd__nand2_1
X_13882_ _18913_/Q _14081_/B _13842_/X _18889_/Q _13881_/X vssd1 vssd1 vccd1 vccd1
+ _13882_/X sky130_fd_sc_hd__a221o_1
XFILLER_189_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15621_ _18144_/Q _15772_/B vssd1 vssd1 vccd1 vccd1 _15736_/A sky130_fd_sc_hd__nand2_2
XTAP_2020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12833_ _12646_/B _12793_/Y _12597_/B _17953_/Q vssd1 vssd1 vccd1 vccd1 _12833_/X
+ sky130_fd_sc_hd__a2bb2o_1
XTAP_2031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_222_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18340_ _18374_/CLK _18340_/D vssd1 vssd1 vccd1 vccd1 _18340_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15552_ _15558_/B _15550_/X _15551_/X _15536_/X vssd1 vssd1 vccd1 vccd1 _18468_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_1330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12764_ _12940_/A vssd1 vssd1 vccd1 vccd1 _12764_/X sky130_fd_sc_hd__buf_4
XTAP_2075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14503_ _14503_/A vssd1 vssd1 vccd1 vccd1 _18225_/D sky130_fd_sc_hd__clkbuf_1
X_11715_ _11683_/X _11697_/X _11705_/X _11598_/B _11714_/X vssd1 vssd1 vccd1 vccd1
+ _11716_/B sky130_fd_sc_hd__a2111o_1
X_15483_ _18487_/Q _18451_/Q _15494_/S vssd1 vssd1 vccd1 vccd1 _15483_/X sky130_fd_sc_hd__mux2_1
XFILLER_163_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18271_ _18275_/CLK _18271_/D vssd1 vssd1 vccd1 vccd1 _18271_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12695_ _12691_/B _12613_/A _12693_/Y _12694_/X _12667_/X vssd1 vssd1 vccd1 vccd1
+ _17935_/D sky130_fd_sc_hd__a221o_1
XTAP_1396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_159_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17222_ _17222_/A vssd1 vssd1 vccd1 vccd1 _17464_/A sky130_fd_sc_hd__buf_2
X_11646_ _17862_/Q vssd1 vssd1 vccd1 vccd1 _12251_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_14434_ _14404_/A _09502_/B _14386_/B vssd1 vssd1 vccd1 vccd1 _14434_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_128_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14365_ _14373_/C _14365_/B vssd1 vssd1 vccd1 vccd1 _14381_/A sky130_fd_sc_hd__nand2_1
X_17153_ _17156_/B _17151_/X _17152_/Y _17140_/X vssd1 vssd1 vccd1 vccd1 _18850_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_128_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11577_ _11577_/A _11577_/B _11549_/X vssd1 vssd1 vccd1 vccd1 _11578_/A sky130_fd_sc_hd__or3b_1
XFILLER_200_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16104_ _16109_/B _16101_/X _16103_/X _16097_/X vssd1 vssd1 vccd1 vccd1 _18600_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_122_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13316_ _18090_/Q _13313_/X _13315_/Y _13074_/X vssd1 vssd1 vccd1 vccd1 _18090_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_183_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17084_ _17148_/A vssd1 vssd1 vccd1 vccd1 _17136_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_10528_ _10899_/A _10528_/B vssd1 vssd1 vccd1 vccd1 _10528_/X sky130_fd_sc_hd__and2_1
XFILLER_128_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14296_ _14296_/A _14296_/B vssd1 vssd1 vccd1 vccd1 _14296_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_6_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16035_ _18622_/Q _18586_/Q _16050_/S vssd1 vssd1 vccd1 vccd1 _16035_/X sky130_fd_sc_hd__mux2_1
XFILLER_182_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13247_ _13255_/A _18078_/Q vssd1 vssd1 vccd1 vccd1 _13248_/A sky130_fd_sc_hd__and2_1
XFILLER_143_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10459_ _10932_/A _10512_/B _10459_/C vssd1 vssd1 vccd1 vccd1 _10459_/X sky130_fd_sc_hd__and3_1
XFILLER_108_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13178_ _13186_/A _18047_/Q vssd1 vssd1 vccd1 vccd1 _13179_/A sky130_fd_sc_hd__and2_1
XFILLER_44_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12129_ _12129_/A vssd1 vssd1 vccd1 vccd1 _13649_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_85_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17986_ _17987_/CLK _17986_/D vssd1 vssd1 vccd1 vccd1 _17986_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_28_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16937_ _16943_/B _16934_/X _16936_/X _16917_/X vssd1 vssd1 vccd1 vccd1 _18798_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_38_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_93_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16868_ _16928_/A vssd1 vssd1 vccd1 vccd1 _16900_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_225_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_203_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18607_ _18607_/CLK _18607_/D vssd1 vssd1 vccd1 vccd1 _18607_/Q sky130_fd_sc_hd__dfxtp_2
X_15819_ _15818_/B _15817_/X _15818_/Y _15803_/X vssd1 vssd1 vccd1 vccd1 _18533_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_20_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_213_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16799_ _16813_/A _16803_/B vssd1 vssd1 vccd1 vccd1 _16799_/Y sky130_fd_sc_hd__nand2_1
XFILLER_129_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09340_ _18434_/Q _18433_/Q _18432_/Q vssd1 vssd1 vccd1 vccd1 _09344_/A sky130_fd_sc_hd__or3_4
X_18538_ _18572_/CLK _18538_/D vssd1 vssd1 vccd1 vccd1 _18538_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_52_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09271_ _09271_/A _09271_/B _09271_/C vssd1 vssd1 vccd1 vccd1 _09440_/A sky130_fd_sc_hd__and3_2
XFILLER_209_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18469_ _18469_/CLK _18469_/D vssd1 vssd1 vccd1 vccd1 _18469_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_21_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_155_wb_clk_i _18102_/CLK vssd1 vssd1 vccd1 vccd1 _18125_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_140_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_228_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_180_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_228_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_216_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08986_ _08998_/A vssd1 vssd1 vccd1 vccd1 _08991_/A sky130_fd_sc_hd__buf_12
XTAP_5629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_228_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_113_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_186_1346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09607_ _10124_/A _13005_/A _09606_/Y vssd1 vssd1 vccd1 vccd1 _09608_/B sky130_fd_sc_hd__a21o_1
XFILLER_83_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_231_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_189_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_188_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09538_ _18114_/Q _09540_/B vssd1 vssd1 vccd1 vccd1 _09589_/B sky130_fd_sc_hd__and2_2
XFILLER_227_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_231_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_212_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09469_ _09475_/A _09463_/X _09466_/B _18138_/D vssd1 vssd1 vccd1 vccd1 _18137_/D
+ sky130_fd_sc_hd__a31o_1
XPHY_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_196_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11500_ _13509_/A _11496_/Y _11455_/D _11499_/X vssd1 vssd1 vccd1 vccd1 _11500_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_12_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12480_ _17907_/Q _12487_/B _12484_/A vssd1 vssd1 vccd1 vccd1 _12480_/Y sky130_fd_sc_hd__a21boi_1
XFILLER_132_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_200_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11431_ _11431_/A _11431_/B vssd1 vssd1 vccd1 vccd1 _11431_/Y sky130_fd_sc_hd__nor2_1
XFILLER_22_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14150_ _14143_/X _14149_/X _12022_/C vssd1 vssd1 vccd1 vccd1 _14150_/X sky130_fd_sc_hd__o21a_1
XFILLER_153_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11362_ _11617_/B _11447_/A vssd1 vssd1 vccd1 vccd1 _11790_/B sky130_fd_sc_hd__nor2_2
XFILLER_165_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19106__77 vssd1 vssd1 vccd1 vccd1 _19106__77/HI _19214_/A sky130_fd_sc_hd__conb_1
XFILLER_137_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13101_ _13107_/A _18012_/Q vssd1 vssd1 vccd1 vccd1 _13102_/A sky130_fd_sc_hd__and2_1
XFILLER_153_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10313_ _12131_/A _12133_/A vssd1 vssd1 vccd1 vccd1 _10313_/Y sky130_fd_sc_hd__nor2_1
XFILLER_180_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14081_ _18482_/Q _14081_/B vssd1 vssd1 vccd1 vccd1 _14081_/X sky130_fd_sc_hd__and2_1
XFILLER_3_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11293_ _17789_/Q _17788_/Q _17790_/Q vssd1 vssd1 vccd1 vccd1 _11951_/B sky130_fd_sc_hd__o21a_2
XFILLER_65_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13032_ _17989_/Q _13036_/B vssd1 vssd1 vccd1 vccd1 _13032_/X sky130_fd_sc_hd__or2_1
Xclkbuf_5_22_0_wb_clk_i clkbuf_5_23_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _18144_/CLK
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_79_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10244_ _10412_/A vssd1 vssd1 vccd1 vccd1 _12032_/A sky130_fd_sc_hd__buf_6
XFILLER_133_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17840_ _17890_/CLK _17840_/D vssd1 vssd1 vccd1 vccd1 _17840_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_65_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10175_ _10175_/A _10175_/B vssd1 vssd1 vccd1 vccd1 _10422_/A sky130_fd_sc_hd__xor2_2
XFILLER_121_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17771_ _19029_/Q _12323_/C _14436_/X vssd1 vssd1 vccd1 vccd1 _19029_/D sky130_fd_sc_hd__o21a_1
XFILLER_78_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14983_ _14995_/A _14983_/B vssd1 vssd1 vccd1 vccd1 _14983_/Y sky130_fd_sc_hd__nand2_1
XFILLER_93_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16722_ _18785_/Q _18749_/Q _16742_/S vssd1 vssd1 vccd1 vccd1 _16722_/X sky130_fd_sc_hd__mux2_1
X_13934_ _18322_/Q _13723_/X _13743_/X _18304_/Q vssd1 vssd1 vccd1 vccd1 _13934_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_75_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16653_ _16658_/B _16651_/X _16652_/X _16639_/X vssd1 vssd1 vccd1 vccd1 _18732_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_170_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13865_ _18814_/Q _13577_/X _13860_/X _13864_/X vssd1 vssd1 vccd1 vccd1 _13865_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_228_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_223_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15604_ _18518_/Q _18482_/Q _15604_/S vssd1 vssd1 vccd1 vccd1 _15604_/X sky130_fd_sc_hd__mux2_1
XFILLER_34_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12816_ _17949_/Q vssd1 vssd1 vccd1 vccd1 _12816_/X sky130_fd_sc_hd__clkbuf_2
X_16584_ _16828_/A vssd1 vssd1 vccd1 vccd1 _16631_/A sky130_fd_sc_hd__clkbuf_2
X_13796_ _18273_/Q _13733_/X _13792_/X _13795_/X vssd1 vssd1 vccd1 vccd1 _13796_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_163_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18323_ _18350_/CLK _18323_/D vssd1 vssd1 vccd1 vccd1 _18323_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_128_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15535_ _15739_/A vssd1 vssd1 vccd1 vccd1 _15616_/A sky130_fd_sc_hd__clkbuf_2
XTAP_1160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12747_ _12748_/B _12747_/B vssd1 vssd1 vccd1 vccd1 _12747_/Y sky130_fd_sc_hd__nand2_1
XFILLER_187_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18254_ _18254_/CLK _18254_/D vssd1 vssd1 vccd1 vccd1 _18254_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_128_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15466_ _16055_/A _15599_/C vssd1 vssd1 vccd1 vccd1 _15473_/B sky130_fd_sc_hd__nor2_2
XFILLER_187_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12678_ _12691_/B _12646_/A _12672_/Y vssd1 vssd1 vccd1 vccd1 _12679_/B sky130_fd_sc_hd__o21ai_1
XFILLER_124_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17205_ _18182_/Q vssd1 vssd1 vccd1 vccd1 _17448_/A sky130_fd_sc_hd__clkbuf_2
X_11629_ _11615_/Y _11624_/X _11603_/B vssd1 vssd1 vccd1 vccd1 _11629_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_8_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14417_ _14420_/A _14417_/B vssd1 vssd1 vccd1 vccd1 _18194_/D sky130_fd_sc_hd__nor2_1
XFILLER_204_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18185_ _18230_/CLK _18185_/D vssd1 vssd1 vccd1 vccd1 _18185_/Q sky130_fd_sc_hd__dfxtp_1
X_15397_ _15423_/A _15997_/B _15423_/C vssd1 vssd1 vccd1 vccd1 _15397_/X sky130_fd_sc_hd__or3_1
XFILLER_200_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17136_ _17136_/A _17425_/B _17173_/C vssd1 vssd1 vccd1 vccd1 _17136_/X sky130_fd_sc_hd__or3_1
XFILLER_184_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14348_ _18181_/Q vssd1 vssd1 vccd1 vccd1 _15607_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_171_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17067_ _18866_/Q _18830_/Q _17074_/S vssd1 vssd1 vccd1 vccd1 _17067_/X sky130_fd_sc_hd__mux2_1
X_14279_ _14279_/A _14323_/B vssd1 vssd1 vccd1 vccd1 _14296_/A sky130_fd_sc_hd__nor2_1
XFILLER_170_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16018_ _16017_/B _16015_/X _16017_/Y _16008_/X vssd1 vssd1 vccd1 vccd1 _18581_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19120__91 vssd1 vssd1 vccd1 vccd1 _19120__91/HI _19228_/A sky130_fd_sc_hd__conb_1
XFILLER_170_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17969_ _17969_/CLK _17969_/D vssd1 vssd1 vccd1 vccd1 _17969_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_100_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_214_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_226_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_230_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_213_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09323_ _18524_/Q _18523_/Q _18522_/Q vssd1 vssd1 vccd1 vccd1 _09327_/A sky130_fd_sc_hd__or3_4
XFILLER_94_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_230_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09254_ _09254_/A _09254_/B _09254_/C vssd1 vssd1 vccd1 vccd1 _09254_/Y sky130_fd_sc_hd__nand3_4
XFILLER_166_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_221_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09185_ _18614_/Q _18613_/Q _18612_/Q vssd1 vssd1 vccd1 vccd1 _09186_/D sky130_fd_sc_hd__or3_4
XFILLER_222_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_218_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_52_wb_clk_i clkbuf_5_16_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18821_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_4725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08969_ _08972_/A vssd1 vssd1 vccd1 vccd1 _08969_/Y sky130_fd_sc_hd__inv_2
XTAP_4736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11980_ _11980_/A _11980_/B _12025_/A _12025_/D vssd1 vssd1 vccd1 vccd1 _12022_/B
+ sky130_fd_sc_hd__and4_1
XTAP_4769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_216_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_205_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10931_ _09304_/B _09294_/D _09294_/A _10569_/A _10542_/X _10518_/X vssd1 vssd1 vccd1
+ vccd1 _10932_/B sky130_fd_sc_hd__mux4_2
XFILLER_17_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_216_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_231_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13650_ _13664_/A vssd1 vssd1 vccd1 vccd1 _13733_/A sky130_fd_sc_hd__buf_6
XFILLER_140_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10862_ _09695_/X _09696_/X _09697_/X _09698_/X _10852_/X _12089_/A vssd1 vssd1 vccd1
+ vccd1 _10862_/X sky130_fd_sc_hd__mux4_2
XFILLER_72_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12601_ _12600_/A _12600_/C _12600_/B vssd1 vssd1 vccd1 vccd1 _12601_/X sky130_fd_sc_hd__a21o_1
XFILLER_169_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13581_ _13702_/A vssd1 vssd1 vccd1 vccd1 _13581_/X sky130_fd_sc_hd__buf_6
XFILLER_140_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10793_ _09209_/A _09219_/B _09214_/D _09214_/B _10770_/X _10695_/A vssd1 vssd1 vccd1
+ vccd1 _10793_/X sky130_fd_sc_hd__mux4_2
XPHY_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_213_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15320_ _15373_/A _15325_/B vssd1 vssd1 vccd1 vccd1 _15320_/Y sky130_fd_sc_hd__nand2_1
X_12532_ _12523_/X _12535_/A _12531_/X _12147_/X vssd1 vssd1 vccd1 vccd1 _17916_/D
+ sky130_fd_sc_hd__o211ai_1
XFILLER_185_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_149_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15251_ _18437_/Q _18401_/Q _15267_/S vssd1 vssd1 vccd1 vccd1 _15251_/X sky130_fd_sc_hd__mux2_1
X_12463_ _17904_/Q _17903_/Q _12487_/B vssd1 vssd1 vccd1 vccd1 _12466_/C sky130_fd_sc_hd__o21ai_1
XFILLER_201_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11414_ _17883_/Q vssd1 vssd1 vccd1 vccd1 _11415_/B sky130_fd_sc_hd__inv_2
X_14202_ _14275_/A vssd1 vssd1 vccd1 vccd1 _14202_/X sky130_fd_sc_hd__clkbuf_2
X_15182_ _15182_/A _15182_/B vssd1 vssd1 vccd1 vccd1 _15182_/Y sky130_fd_sc_hd__nand2_1
XFILLER_201_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12394_ _17896_/Q _12394_/B _12394_/C vssd1 vssd1 vccd1 vccd1 _12395_/B sky130_fd_sc_hd__nor3_1
XFILLER_32_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14133_ _18299_/Q _13940_/X _14131_/X _14132_/X vssd1 vssd1 vccd1 vccd1 _14133_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_137_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11345_ _11345_/A _11385_/A vssd1 vssd1 vccd1 vccd1 _11388_/A sky130_fd_sc_hd__nor2_1
XFILLER_67_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_153_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14064_ _18410_/Q _13612_/A _14027_/A _18401_/Q _14063_/X vssd1 vssd1 vccd1 vccd1
+ _14064_/X sky130_fd_sc_hd__a221o_4
XFILLER_3_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18941_ _18965_/CLK _18941_/D vssd1 vssd1 vccd1 vccd1 _18941_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_153_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11276_ _11282_/B _11832_/B _11275_/X _11807_/A vssd1 vssd1 vccd1 vccd1 _11277_/C
+ sky130_fd_sc_hd__o22a_1
XFILLER_4_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_152_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13015_ _13025_/A vssd1 vssd1 vccd1 vccd1 _13015_/X sky130_fd_sc_hd__clkbuf_2
X_10227_ _10440_/A _10227_/B vssd1 vssd1 vccd1 vccd1 _10560_/S sky130_fd_sc_hd__xnor2_4
X_18872_ _18875_/CLK _18872_/D vssd1 vssd1 vccd1 vccd1 _18872_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_121_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17823_ _17824_/CLK _17823_/D vssd1 vssd1 vccd1 vccd1 _17823_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10158_ _10158_/A _10165_/S vssd1 vssd1 vccd1 vccd1 _10159_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3 hold3/A vssd1 vssd1 vccd1 vccd1 hold3/X sky130_fd_sc_hd__clkdlybuf4s50_1
XTAP_5971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17754_ _17756_/A _19021_/Q vssd1 vssd1 vccd1 vccd1 _17755_/A sky130_fd_sc_hd__and2_1
XFILLER_66_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_181_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14966_ _14971_/B _14964_/X _14965_/X _14961_/X vssd1 vssd1 vccd1 vccd1 _18330_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_43_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10089_ _09248_/B _09243_/B _10089_/S vssd1 vssd1 vccd1 vccd1 _10089_/X sky130_fd_sc_hd__mux2_1
XFILLER_48_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_1330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16705_ _16712_/B _16702_/X _16703_/X _16704_/X vssd1 vssd1 vccd1 vccd1 _18744_/D
+ sky130_fd_sc_hd__o211a_1
X_13917_ _18739_/Q _13642_/X _13841_/A _18745_/Q vssd1 vssd1 vccd1 vccd1 _13917_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_47_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17685_ _17712_/A _17685_/B vssd1 vssd1 vccd1 vccd1 _17686_/A sky130_fd_sc_hd__and2_1
X_14897_ _14932_/A _14900_/B vssd1 vssd1 vccd1 vccd1 _14897_/Y sky130_fd_sc_hd__nand2_1
XFILLER_130_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_223_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16636_ _16783_/A _16650_/B vssd1 vssd1 vccd1 vccd1 _16648_/B sky130_fd_sc_hd__nor2_2
XFILLER_23_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13848_ _13848_/A vssd1 vssd1 vccd1 vccd1 _13848_/X sky130_fd_sc_hd__buf_6
XFILLER_74_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16567_ _16808_/A vssd1 vssd1 vccd1 vccd1 _16615_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_22_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13779_ _18660_/Q _13714_/X _13698_/A _18651_/Q _13778_/X vssd1 vssd1 vccd1 vccd1
+ _13779_/X sky130_fd_sc_hd__a221o_2
XFILLER_95_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_203_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18306_ _18308_/CLK _18306_/D vssd1 vssd1 vccd1 vccd1 _18306_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_31_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15518_ _15568_/A vssd1 vssd1 vccd1 vccd1 _15545_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_176_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_203_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16498_ _18731_/Q _18695_/Q _16509_/S vssd1 vssd1 vccd1 vccd1 _16498_/X sky130_fd_sc_hd__mux2_1
XFILLER_31_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18237_ _18263_/CLK _18237_/D vssd1 vssd1 vccd1 vccd1 _18237_/Q sky130_fd_sc_hd__dfxtp_1
X_15449_ _18480_/Q _18444_/Q _15458_/S vssd1 vssd1 vccd1 vccd1 _15449_/X sky130_fd_sc_hd__mux2_1
XFILLER_175_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18168_ _18182_/CLK _18168_/D vssd1 vssd1 vccd1 vccd1 _18168_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_11_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17119_ _17119_/A _17119_/B _18178_/Q _18177_/Q vssd1 vssd1 vccd1 vccd1 _17549_/B
+ sky130_fd_sc_hd__or4_4
XFILLER_102_1277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18099_ _18110_/CLK _18099_/D vssd1 vssd1 vccd1 vccd1 _18099_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_102_1299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09941_ _09936_/X _09938_/X _10305_/S vssd1 vssd1 vccd1 vccd1 _09941_/X sky130_fd_sc_hd__mux2_1
X_19097__68 vssd1 vssd1 vccd1 vccd1 _19097__68/HI _19205_/A sky130_fd_sc_hd__conb_1
XFILLER_48_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09872_ _09872_/A _09872_/B vssd1 vssd1 vccd1 vccd1 _09872_/Y sky130_fd_sc_hd__nor2_1
XTAP_741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_219_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_225_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_218_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINSDIODE2_16 _09209_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_27 _09458_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_38 _09937_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_1306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINSDIODE2_49 _10528_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_227_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_214_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_213_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_170_wb_clk_i clkbuf_5_11_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18052_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_09306_ _18449_/Q _18448_/Q _18447_/Q vssd1 vssd1 vccd1 vccd1 _10575_/A sky130_fd_sc_hd__or3_4
XFILLER_16_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09237_ _09237_/A _09237_/B _09237_/C _09237_/D vssd1 vssd1 vccd1 vccd1 _09238_/C
+ sky130_fd_sc_hd__and4_1
XFILLER_186_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_222_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_1311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09168_ _18659_/Q _18658_/Q _18657_/Q vssd1 vssd1 vccd1 vccd1 _09170_/C sky130_fd_sc_hd__or3_4
XFILLER_166_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_148_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09099_ _18782_/Q _18781_/Q _18780_/Q vssd1 vssd1 vccd1 vccd1 _09103_/A sky130_fd_sc_hd__or3_4
XFILLER_163_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11130_ _17800_/Q vssd1 vssd1 vccd1 vccd1 _11541_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_218_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11061_ _11336_/A vssd1 vssd1 vccd1 vccd1 _13427_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_62_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_231_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10012_ _10001_/X _10011_/X _09657_/X vssd1 vssd1 vccd1 vccd1 _10012_/X sky130_fd_sc_hd__o21a_1
XFILLER_118_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14820_ _14827_/B _14817_/X _14818_/X _14819_/X vssd1 vssd1 vccd1 vccd1 _18294_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_76_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14751_ _14753_/B _14749_/X _14750_/Y _14738_/X vssd1 vssd1 vccd1 vccd1 _18277_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_229_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_217_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11963_ _11963_/A _11985_/A vssd1 vssd1 vccd1 vccd1 _12026_/D sky130_fd_sc_hd__nor2_1
XTAP_3865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13702_ _13702_/A vssd1 vssd1 vccd1 vccd1 _13834_/A sky130_fd_sc_hd__buf_4
XTAP_3887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17470_ _17469_/B _17467_/X _17469_/Y _17461_/X vssd1 vssd1 vccd1 vccd1 _18929_/D
+ sky130_fd_sc_hd__o211a_1
X_10914_ _11925_/A _10914_/B vssd1 vssd1 vccd1 vccd1 _10914_/X sky130_fd_sc_hd__and2_1
XFILLER_229_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14682_ _18262_/Q _14683_/B _14681_/Y _14668_/X vssd1 vssd1 vccd1 vccd1 _18262_/D
+ sky130_fd_sc_hd__o211a_1
X_11894_ _09069_/B _11879_/A _11893_/Y vssd1 vssd1 vccd1 vccd1 _17837_/D sky130_fd_sc_hd__a21o_1
XFILLER_44_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_189_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16421_ _18711_/Q _18675_/Q _16421_/S vssd1 vssd1 vccd1 vccd1 _16421_/X sky130_fd_sc_hd__mux2_1
XFILLER_72_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13633_ _18465_/Q _13525_/A _13621_/X _18468_/Q _13632_/X vssd1 vssd1 vccd1 vccd1
+ _13633_/X sky130_fd_sc_hd__a221o_1
X_10845_ _09126_/C _09131_/B _09136_/D _09131_/D _10882_/S _10824_/A vssd1 vssd1 vccd1
+ vccd1 _10845_/X sky130_fd_sc_hd__mux4_2
XFILLER_38_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19140_ _19140_/A _09034_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[10] sky130_fd_sc_hd__ebufn_8
XFILLER_213_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16352_ _18695_/Q _18659_/Q _16363_/S vssd1 vssd1 vccd1 vccd1 _16352_/X sky130_fd_sc_hd__mux2_1
XFILLER_198_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13564_ _13772_/A vssd1 vssd1 vccd1 vccd1 _13715_/A sky130_fd_sc_hd__buf_4
XFILLER_125_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10776_ _09294_/C _09299_/B _09304_/D _09299_/D _10716_/A _10701_/A vssd1 vssd1 vccd1
+ vccd1 _10777_/B sky130_fd_sc_hd__mux4_1
XFILLER_12_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15303_ _15303_/A _15303_/B vssd1 vssd1 vccd1 vccd1 _15303_/Y sky130_fd_sc_hd__nand2_1
XFILLER_9_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_200_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12515_ _12521_/A vssd1 vssd1 vccd1 vccd1 _17543_/S sky130_fd_sc_hd__buf_4
X_16283_ _17228_/A vssd1 vssd1 vccd1 vccd1 _16524_/A sky130_fd_sc_hd__buf_2
XFILLER_157_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13495_ _13557_/A _13563_/B vssd1 vssd1 vccd1 vccd1 _13720_/A sky130_fd_sc_hd__nor2_2
XFILLER_8_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18022_ _18095_/CLK _18022_/D vssd1 vssd1 vccd1 vccd1 _18022_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_9_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15234_ _15239_/B _15231_/X _15233_/X _15224_/X vssd1 vssd1 vccd1 vccd1 _18396_/D
+ sky130_fd_sc_hd__o211a_1
X_12446_ _12446_/A _12470_/B vssd1 vssd1 vccd1 vccd1 _12452_/A sky130_fd_sc_hd__or2_1
XFILLER_139_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15165_ _15178_/A _15169_/B vssd1 vssd1 vccd1 vccd1 _15165_/Y sky130_fd_sc_hd__nand2_1
XFILLER_158_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12377_ _12388_/A _12388_/B vssd1 vssd1 vccd1 vccd1 _12379_/B sky130_fd_sc_hd__or2b_1
XFILLER_99_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11328_ _11328_/A _11339_/D vssd1 vssd1 vccd1 vccd1 _11385_/B sky130_fd_sc_hd__nor2_1
X_14116_ _18941_/Q _13532_/A _13539_/A _18917_/Q vssd1 vssd1 vccd1 vccd1 _14116_/X
+ sky130_fd_sc_hd__a22o_1
X_15096_ _15241_/A _15134_/B vssd1 vssd1 vccd1 vccd1 _15107_/B sky130_fd_sc_hd__nor2_2
XFILLER_153_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18924_ _18926_/CLK _18924_/D vssd1 vssd1 vccd1 vccd1 _18924_/Q sky130_fd_sc_hd__dfxtp_4
X_14047_ _18536_/Q _13834_/A _14045_/X _14046_/X vssd1 vssd1 vccd1 vccd1 _14047_/X
+ sky130_fd_sc_hd__a211o_1
X_11259_ _11748_/C _11586_/D vssd1 vssd1 vccd1 vccd1 _11259_/Y sky130_fd_sc_hd__nor2_1
XFILLER_171_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_1362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18855_ _18862_/CLK _18855_/D vssd1 vssd1 vccd1 vccd1 _18855_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_67_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_227_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17806_ _17806_/CLK _17806_/D vssd1 vssd1 vccd1 vccd1 _17806_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_10_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18786_ _18786_/CLK _18786_/D vssd1 vssd1 vccd1 vccd1 _18786_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_227_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15998_ _16003_/B _15995_/X _15997_/X _15988_/X vssd1 vssd1 vccd1 vccd1 _18576_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_94_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17737_ _17745_/A _19013_/Q vssd1 vssd1 vccd1 vccd1 _17738_/A sky130_fd_sc_hd__and2_1
XFILLER_78_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14949_ _14995_/A _14949_/B vssd1 vssd1 vccd1 vccd1 _14949_/Y sky130_fd_sc_hd__nand2_1
XFILLER_36_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17668_ _17641_/X _17663_/Y _17654_/X _17664_/Y _18979_/Q vssd1 vssd1 vccd1 vccd1
+ _17669_/B sky130_fd_sc_hd__a32o_1
XINSDIODE2_120 _15233_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINSDIODE2_131 _16431_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_142 _17265_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_153 _18422_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16619_ _16659_/A vssd1 vssd1 vccd1 vccd1 _16619_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_126_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_211_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XINSDIODE2_164 _18361_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17599_ _17571_/X _17590_/Y _17582_/X _17592_/Y _18962_/Q vssd1 vssd1 vccd1 vccd1
+ _17600_/B sky130_fd_sc_hd__a32o_1
XINSDIODE2_175 _18712_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_186 _09098_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_206_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_197 _10518_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_1333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09022_ _09022_/A vssd1 vssd1 vccd1 vccd1 _09022_/Y sky130_fd_sc_hd__inv_2
XFILLER_108_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_4_3_0_wb_clk_i clkbuf_4_3_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_5_7_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_145_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09924_ _09924_/A vssd1 vssd1 vccd1 vccd1 _10376_/B sky130_fd_sc_hd__buf_2
XFILLER_217_1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09855_ _09855_/A _09855_/B vssd1 vssd1 vccd1 vccd1 _09858_/A sky130_fd_sc_hd__xor2_4
XFILLER_24_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_150_1348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09786_ _10213_/A _09780_/B _09785_/X vssd1 vssd1 vccd1 vccd1 _09787_/B sky130_fd_sc_hd__o21a_1
XFILLER_86_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_227_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_199_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_1282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_230_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_215_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_197_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10630_ _10625_/B _12958_/A vssd1 vssd1 vccd1 vccd1 _10630_/X sky130_fd_sc_hd__and2b_1
XFILLER_198_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_201_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_210_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10561_ _10559_/X _10560_/X _10561_/S vssd1 vssd1 vccd1 vccd1 _10561_/X sky130_fd_sc_hd__mux2_1
XFILLER_10_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12300_ _12300_/A _12300_/B vssd1 vssd1 vccd1 vccd1 _12301_/A sky130_fd_sc_hd__and2_1
X_13280_ _19002_/Q _19001_/Q _19004_/Q _19003_/Q vssd1 vssd1 vccd1 vccd1 _13281_/B
+ sky130_fd_sc_hd__or4_1
XFILLER_212_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10492_ _10454_/X _10489_/X _10491_/X _10923_/S vssd1 vssd1 vccd1 vccd1 _10492_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_154_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12231_ _12231_/A vssd1 vssd1 vccd1 vccd1 _17856_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_108_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_107_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12162_ _12940_/A vssd1 vssd1 vccd1 vccd1 _14436_/A sky130_fd_sc_hd__buf_2
XFILLER_163_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11113_ _13447_/A _11181_/A _11113_/S vssd1 vssd1 vccd1 vccd1 _11114_/A sky130_fd_sc_hd__mux2_1
XFILLER_151_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16970_ _18842_/Q _18806_/Q _16970_/S vssd1 vssd1 vccd1 vccd1 _16970_/X sky130_fd_sc_hd__mux2_1
X_12093_ _14247_/A _13509_/B _12091_/X _12092_/Y vssd1 vssd1 vccd1 vccd1 _12095_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_96_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15921_ _15921_/A _15921_/B _15964_/C vssd1 vssd1 vccd1 vccd1 _15921_/X sky130_fd_sc_hd__or3_1
XTAP_5020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11044_ _11044_/A _11044_/B vssd1 vssd1 vccd1 vccd1 _13346_/A sky130_fd_sc_hd__nand2_1
XFILLER_7_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18640_ _18641_/CLK _18640_/D vssd1 vssd1 vccd1 vccd1 _18640_/Q sky130_fd_sc_hd__dfxtp_4
XTAP_5064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15852_ _18578_/Q _18542_/Q _15859_/S vssd1 vssd1 vccd1 vccd1 _15852_/X sky130_fd_sc_hd__mux2_1
XTAP_5075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14803_ _14802_/B _14801_/X _14802_/Y _14799_/X vssd1 vssd1 vccd1 vccd1 _18290_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_18_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18571_ _18571_/CLK _18571_/D vssd1 vssd1 vccd1 vccd1 _18571_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_4374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_218_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15783_ _15823_/A vssd1 vssd1 vccd1 vccd1 _15783_/X sky130_fd_sc_hd__clkbuf_2
XTAP_4385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12995_ _12990_/Y _12775_/A _12989_/A vssd1 vssd1 vccd1 vccd1 _12995_/X sky130_fd_sc_hd__a21o_1
XFILLER_92_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17522_ _17524_/B _17520_/X _17521_/Y _17517_/X vssd1 vssd1 vccd1 vccd1 _18943_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_3673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14734_ _14734_/A _15175_/B _14757_/C vssd1 vssd1 vccd1 vccd1 _14734_/X sky130_fd_sc_hd__or3_1
XFILLER_17_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11946_ _11964_/C vssd1 vssd1 vccd1 vccd1 _11946_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_75_1216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_205_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_229_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17453_ _17453_/A _17456_/B vssd1 vssd1 vccd1 vccd1 _17453_/Y sky130_fd_sc_hd__nand2_1
XFILLER_229_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14665_ _14665_/A _14665_/B _15257_/B vssd1 vssd1 vccd1 vccd1 _14665_/X sky130_fd_sc_hd__or3_1
XFILLER_33_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11877_ _11879_/A _11877_/B vssd1 vssd1 vccd1 vccd1 _17831_/D sky130_fd_sc_hd__nor2_1
XTAP_2994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16404_ _16473_/A vssd1 vssd1 vccd1 vccd1 _16421_/S sky130_fd_sc_hd__clkbuf_2
X_13616_ _13616_/A vssd1 vssd1 vccd1 vccd1 _13617_/A sky130_fd_sc_hd__buf_6
X_17384_ _17383_/B _17382_/X _17383_/Y _17380_/X vssd1 vssd1 vccd1 vccd1 _18908_/D
+ sky130_fd_sc_hd__o211a_1
X_10828_ _12092_/A _10825_/X _10827_/X _10766_/A vssd1 vssd1 vccd1 vccd1 _10828_/X
+ sky130_fd_sc_hd__a211o_1
X_14596_ _18182_/Q vssd1 vssd1 vccd1 vccd1 _14597_/A sky130_fd_sc_hd__buf_2
XFILLER_38_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16335_ _16342_/B _16332_/X _16333_/X _16334_/X vssd1 vssd1 vccd1 vccd1 _18654_/D
+ sky130_fd_sc_hd__o211a_1
X_13547_ _13563_/A _13547_/B vssd1 vssd1 vccd1 vccd1 _13613_/A sky130_fd_sc_hd__nor2_4
XFILLER_9_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10759_ _09314_/B _09319_/A _09319_/C _09309_/C _10858_/S _10738_/A vssd1 vssd1 vccd1
+ vccd1 _10759_/X sky130_fd_sc_hd__mux4_2
XFILLER_186_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_187_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16266_ _16268_/B _16264_/X _16265_/Y _16252_/X vssd1 vssd1 vccd1 vccd1 _18637_/D
+ sky130_fd_sc_hd__o211a_1
X_13478_ _13480_/A _13478_/B vssd1 vssd1 vccd1 vccd1 _18162_/D sky130_fd_sc_hd__nor2_1
XFILLER_145_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18005_ _18213_/CLK _18005_/D vssd1 vssd1 vccd1 vccd1 _18005_/Q sky130_fd_sc_hd__dfxtp_1
X_15217_ _18392_/Q _15216_/B _15216_/Y _15208_/X vssd1 vssd1 vccd1 vccd1 _18392_/D
+ sky130_fd_sc_hd__o211a_1
X_12429_ _12429_/A _12439_/B vssd1 vssd1 vccd1 vccd1 _12430_/C sky130_fd_sc_hd__nand2_1
X_16197_ _16197_/A vssd1 vssd1 vccd1 vccd1 _16215_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_126_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15148_ _15211_/A vssd1 vssd1 vccd1 vccd1 _15277_/B sky130_fd_sc_hd__buf_2
XFILLER_5_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_153_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19067__38 vssd1 vssd1 vccd1 vccd1 _19067__38/HI _19161_/A sky130_fd_sc_hd__conb_1
X_15079_ _15115_/A _15082_/B vssd1 vssd1 vccd1 vccd1 _15079_/Y sky130_fd_sc_hd__nand2_1
XFILLER_141_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18907_ _18907_/CLK _18907_/D vssd1 vssd1 vccd1 vccd1 _18907_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_101_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_206_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_132_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09640_ _09668_/A _09640_/B vssd1 vssd1 vccd1 vccd1 _09653_/A sky130_fd_sc_hd__xnor2_4
X_18838_ _18875_/CLK _18838_/D vssd1 vssd1 vccd1 vccd1 _18838_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_28_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_109_wb_clk_i clkbuf_5_29_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18533_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_49_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09571_ _09600_/A _09569_/X _09570_/X vssd1 vssd1 vccd1 vccd1 _09573_/B sky130_fd_sc_hd__o21ai_1
X_18769_ _18773_/CLK _18769_/D vssd1 vssd1 vccd1 vccd1 _18769_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_71_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_208_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_180_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_208_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_212_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_220_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09005_ _09029_/A vssd1 vssd1 vccd1 vccd1 _09010_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_191_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_219_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_192_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_151_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_219_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_219_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09907_ _09907_/A _09907_/B vssd1 vssd1 vccd1 vccd1 _10348_/A sky130_fd_sc_hd__nand2_4
XFILLER_99_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_219_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_219_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_219_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09838_ _09828_/B _10193_/B _09837_/Y vssd1 vssd1 vccd1 vccd1 _09840_/B sky130_fd_sc_hd__a21bo_2
XFILLER_98_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_219_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19081__52 vssd1 vssd1 vccd1 vccd1 _19081__52/HI _19189_/A sky130_fd_sc_hd__conb_1
XFILLER_6_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09769_ _18110_/Q vssd1 vssd1 vccd1 vccd1 _09777_/A sky130_fd_sc_hd__inv_2
XTAP_2202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11800_ _11781_/Y _11783_/Y _11780_/Y _11781_/A _11799_/X vssd1 vssd1 vccd1 vccd1
+ _11800_/X sky130_fd_sc_hd__o221a_1
XFILLER_55_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12780_ _13085_/A _13082_/A vssd1 vssd1 vccd1 vccd1 _12784_/B sky130_fd_sc_hd__nor2_1
XFILLER_73_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11731_ _17913_/Q _17912_/Q vssd1 vssd1 vccd1 vccd1 _11732_/B sky130_fd_sc_hd__xnor2_4
XTAP_2279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_202_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14450_ _14414_/A _14445_/Y _14386_/B vssd1 vssd1 vccd1 vccd1 _14450_/Y sky130_fd_sc_hd__o21bai_1
X_11662_ _11748_/C _11586_/C _11669_/B vssd1 vssd1 vccd1 vccd1 _11663_/B sky130_fd_sc_hd__a21oi_1
XTAP_1589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13401_ _13405_/B _13401_/B vssd1 vssd1 vccd1 vccd1 _13402_/A sky130_fd_sc_hd__and2_1
X_10613_ _10612_/A _10612_/B _18121_/Q vssd1 vssd1 vccd1 vccd1 _10614_/B sky130_fd_sc_hd__o21ba_1
X_11593_ _11593_/A _11593_/B vssd1 vssd1 vccd1 vccd1 _11593_/Y sky130_fd_sc_hd__nor2_1
X_14381_ _14381_/A _14381_/B vssd1 vssd1 vccd1 vccd1 _14381_/X sky130_fd_sc_hd__or2_1
XFILLER_70_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_168_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_1274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16120_ _16139_/A vssd1 vssd1 vccd1 vccd1 _16120_/X sky130_fd_sc_hd__clkbuf_2
X_13332_ _18095_/Q _12729_/B _12919_/X vssd1 vssd1 vccd1 vccd1 _13332_/Y sky130_fd_sc_hd__a21oi_1
X_10544_ _09386_/D _09381_/D _09376_/C _09381_/B _10518_/A _10542_/X vssd1 vssd1 vccd1
+ vccd1 _10544_/X sky130_fd_sc_hd__mux4_1
XFILLER_128_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_157_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16051_ _16064_/A _16051_/B vssd1 vssd1 vccd1 vccd1 _16051_/Y sky130_fd_sc_hd__nand2_1
XFILLER_183_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13263_ _13263_/A vssd1 vssd1 vccd1 vccd1 _18084_/D sky130_fd_sc_hd__clkbuf_1
X_10475_ _10475_/A vssd1 vssd1 vccd1 vccd1 _10935_/S sky130_fd_sc_hd__buf_4
XFILLER_182_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15002_ _15042_/A _15150_/B _15054_/C vssd1 vssd1 vccd1 vccd1 _15002_/X sky130_fd_sc_hd__or3_1
XFILLER_124_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_182_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12214_ _11704_/A _11706_/A _12205_/A _11685_/X vssd1 vssd1 vccd1 vccd1 _12215_/C
+ sky130_fd_sc_hd__a31o_1
XFILLER_136_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_135_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13194_ _13194_/A vssd1 vssd1 vccd1 vccd1 _18053_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_135_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12145_ _12145_/A vssd1 vssd1 vccd1 vccd1 _12169_/B sky130_fd_sc_hd__dlymetal6s2s_1
Xclkbuf_leaf_7_wb_clk_i _17929_/CLK vssd1 vssd1 vccd1 vccd1 _17931_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_151_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16953_ _18838_/Q _18802_/Q _16970_/S vssd1 vssd1 vccd1 vccd1 _16953_/X sky130_fd_sc_hd__mux2_1
X_12076_ _10218_/A _12975_/A _12075_/Y vssd1 vssd1 vccd1 vccd1 _12077_/B sky130_fd_sc_hd__a21o_1
XFILLER_150_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15904_ _17120_/A _16366_/B vssd1 vssd1 vccd1 vccd1 _15975_/A sky130_fd_sc_hd__or2_1
X_11027_ _11021_/X _09828_/B _11023_/X _11026_/X vssd1 vssd1 vccd1 vccd1 _17781_/D
+ sky130_fd_sc_hd__o211a_1
X_16884_ _16884_/A _16884_/B vssd1 vssd1 vccd1 vccd1 _16884_/Y sky130_fd_sc_hd__nand2_1
Xclkbuf_leaf_202_wb_clk_i clkbuf_5_7_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18953_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_18623_ _18623_/CLK _18623_/D vssd1 vssd1 vccd1 vccd1 _18623_/Q sky130_fd_sc_hd__dfxtp_1
X_15835_ _18574_/Q _18538_/Q _15838_/S vssd1 vssd1 vccd1 vccd1 _15835_/X sky130_fd_sc_hd__mux2_1
XTAP_4160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_225_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18554_ _18557_/CLK _18554_/D vssd1 vssd1 vccd1 vccd1 _18554_/Q sky130_fd_sc_hd__dfxtp_1
X_15766_ _15815_/A _15769_/B vssd1 vssd1 vccd1 vccd1 _15766_/Y sky130_fd_sc_hd__nand2_1
XTAP_3470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12978_ _17986_/Q _12955_/X _12976_/X _12977_/Y _12949_/Y vssd1 vssd1 vccd1 vccd1
+ _12978_/X sky130_fd_sc_hd__a221o_1
XTAP_3481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17505_ _17575_/A vssd1 vssd1 vccd1 vccd1 _17538_/A sky130_fd_sc_hd__clkbuf_2
X_14717_ _18269_/Q _14715_/B _14715_/Y _14716_/X vssd1 vssd1 vccd1 vccd1 _18269_/D
+ sky130_fd_sc_hd__o211a_1
X_18485_ _18485_/CLK _18485_/D vssd1 vssd1 vccd1 vccd1 _18485_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_45_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11929_ _11945_/A _11945_/B vssd1 vssd1 vccd1 vccd1 _11929_/X sky130_fd_sc_hd__and2_1
X_15697_ _15717_/A vssd1 vssd1 vccd1 vccd1 _15714_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_61_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17436_ _18957_/Q _18921_/Q _17447_/S vssd1 vssd1 vccd1 vccd1 _17436_/X sky130_fd_sc_hd__mux2_1
XFILLER_220_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14648_ _18254_/Q _14646_/B _14646_/Y _14647_/X vssd1 vssd1 vccd1 vccd1 _18254_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_221_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_159_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_207_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_159_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_220_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17367_ _18940_/Q _18904_/Q _17367_/S vssd1 vssd1 vccd1 vccd1 _17367_/X sky130_fd_sc_hd__mux2_1
XFILLER_174_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14579_ _17635_/A _17687_/B vssd1 vssd1 vccd1 vccd1 _16850_/A sky130_fd_sc_hd__or2_4
XFILLER_203_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16318_ _16317_/B _16316_/X _16317_/Y _16314_/X vssd1 vssd1 vccd1 vccd1 _18650_/D
+ sky130_fd_sc_hd__o211a_1
X_17298_ _18922_/Q _18886_/Q _17298_/S vssd1 vssd1 vccd1 vccd1 _17298_/X sky130_fd_sc_hd__mux2_1
X_16249_ _16256_/B _16247_/X _16248_/X _16230_/X vssd1 vssd1 vccd1 vccd1 _18633_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_133_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_228_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_228_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_214_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09623_ _09645_/A _09623_/B vssd1 vssd1 vccd1 vccd1 _09665_/A sky130_fd_sc_hd__xnor2_2
XFILLER_23_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09554_ _09568_/A _09537_/B _09553_/Y vssd1 vssd1 vccd1 vccd1 _09555_/B sky130_fd_sc_hd__o21a_1
XFILLER_55_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_1282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_224_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_212_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_224_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09485_ input2/X vssd1 vssd1 vccd1 vccd1 _12224_/A sky130_fd_sc_hd__inv_2
XFILLER_212_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_77_wb_clk_i clkbuf_5_23_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18635_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_197_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_177_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_221_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_192_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_1351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10260_ _11916_/A _11916_/B vssd1 vssd1 vccd1 vccd1 _11910_/B sky130_fd_sc_hd__xnor2_1
XFILLER_156_1310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_5_12_0_wb_clk_i clkbuf_4_6_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_5_12_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_191_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_180_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_1354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10191_ _10191_/A _10258_/B vssd1 vssd1 vccd1 vccd1 _10192_/B sky130_fd_sc_hd__xor2_1
XFILLER_191_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13950_ _18487_/Q _13735_/X _13721_/X _18511_/Q vssd1 vssd1 vccd1 vccd1 _13950_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_4_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12901_ _12904_/C _12901_/B vssd1 vssd1 vccd1 vccd1 _17963_/D sky130_fd_sc_hd__nor2_1
XFILLER_86_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13881_ _18895_/Q _13877_/X _13879_/X _13880_/X vssd1 vssd1 vccd1 vccd1 _13881_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_100_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_219_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15620_ _15915_/A _15748_/C vssd1 vssd1 vccd1 vccd1 _15633_/B sky130_fd_sc_hd__nor2_1
XFILLER_189_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12832_ _17965_/Q vssd1 vssd1 vccd1 vccd1 _12832_/Y sky130_fd_sc_hd__inv_2
XFILLER_34_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15551_ _15551_/A _15997_/B _15574_/C vssd1 vssd1 vccd1 vccd1 _15551_/X sky130_fd_sc_hd__or3_1
XTAP_1320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12763_ _17940_/Q vssd1 vssd1 vccd1 vccd1 _14373_/A sky130_fd_sc_hd__buf_2
XFILLER_61_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14502_ _18225_/Q _14502_/B vssd1 vssd1 vccd1 vccd1 _14503_/A sky130_fd_sc_hd__and2_1
XTAP_1353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18270_ _18275_/CLK _18270_/D vssd1 vssd1 vccd1 vccd1 _18270_/Q sky130_fd_sc_hd__dfxtp_1
X_11714_ _11711_/X _11714_/B vssd1 vssd1 vccd1 vccd1 _11714_/X sky130_fd_sc_hd__and2b_1
XTAP_1364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15482_ _15487_/B _15480_/X _15481_/X _15474_/X vssd1 vssd1 vccd1 vccd1 _18450_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_203_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_202_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12694_ _12693_/A _12693_/B _12537_/S vssd1 vssd1 vccd1 vccd1 _12694_/X sky130_fd_sc_hd__o21a_1
XFILLER_226_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17221_ _18904_/Q _18868_/Q _17221_/S vssd1 vssd1 vccd1 vccd1 _17221_/X sky130_fd_sc_hd__mux2_1
XFILLER_35_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14433_ _14452_/A _14433_/B vssd1 vssd1 vccd1 vccd1 _18198_/D sky130_fd_sc_hd__nor2_1
X_11645_ _11645_/A _11673_/A vssd1 vssd1 vccd1 vccd1 _11645_/X sky130_fd_sc_hd__or2_1
XFILLER_30_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_1366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17152_ _17152_/A _17156_/B vssd1 vssd1 vccd1 vccd1 _17152_/Y sky130_fd_sc_hd__nand2_1
X_14364_ _14383_/C _18131_/Q _16673_/A vssd1 vssd1 vccd1 vccd1 _14365_/B sky130_fd_sc_hd__or3b_2
XFILLER_168_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11576_ _11556_/X _11701_/A _11575_/X _11563_/B vssd1 vssd1 vccd1 vccd1 _11577_/A
+ sky130_fd_sc_hd__o22a_1
X_16103_ _16115_/A _16703_/B _16115_/C vssd1 vssd1 vccd1 vccd1 _16103_/X sky130_fd_sc_hd__or3_1
XFILLER_183_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13315_ _18090_/Q _13310_/A _13324_/A vssd1 vssd1 vccd1 vccd1 _13315_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_143_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10527_ _09165_/D _09170_/C _09170_/A _09160_/D _10429_/X _10430_/X vssd1 vssd1 vccd1
+ vccd1 _10528_/B sky130_fd_sc_hd__mux4_2
XFILLER_128_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17083_ _18870_/Q _18834_/Q _17094_/S vssd1 vssd1 vccd1 vccd1 _17083_/X sky130_fd_sc_hd__mux2_1
XFILLER_122_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14295_ _14295_/A _14233_/A vssd1 vssd1 vccd1 vccd1 _14296_/B sky130_fd_sc_hd__or2b_1
XFILLER_109_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16034_ _16034_/A vssd1 vssd1 vccd1 vccd1 _16050_/S sky130_fd_sc_hd__clkbuf_2
X_13246_ _13257_/A vssd1 vssd1 vccd1 vccd1 _13255_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_100_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10458_ _09237_/B _09227_/D _09227_/A _10826_/A _10484_/A _10489_/S vssd1 vssd1 vccd1
+ vccd1 _10459_/C sky130_fd_sc_hd__mux4_1
XFILLER_170_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10389_ _10389_/A _10391_/B vssd1 vssd1 vccd1 vccd1 _10389_/X sky130_fd_sc_hd__or2_1
X_13177_ _13199_/A vssd1 vssd1 vccd1 vccd1 _13186_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_112_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12128_ _12128_/A _13494_/B vssd1 vssd1 vccd1 vccd1 _12132_/B sky130_fd_sc_hd__xnor2_1
XFILLER_2_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17985_ _18044_/CLK _17985_/D vssd1 vssd1 vccd1 vccd1 _17985_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16936_ _16936_/A _17516_/B _16936_/C vssd1 vssd1 vccd1 vccd1 _16936_/X sky130_fd_sc_hd__or3_1
XFILLER_133_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12059_ _12059_/A _12089_/B vssd1 vssd1 vccd1 vccd1 _12059_/Y sky130_fd_sc_hd__nand2_1
XFILLER_42_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_211_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16867_ _16874_/B _16864_/X _16866_/X _16848_/X vssd1 vssd1 vccd1 vccd1 _18783_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_37_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15818_ _15818_/A _15818_/B vssd1 vssd1 vccd1 vccd1 _15818_/Y sky130_fd_sc_hd__nand2_1
X_18606_ _18607_/CLK _18606_/D vssd1 vssd1 vccd1 vccd1 _18606_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_80_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16798_ _18805_/Q _18769_/Q _16802_/S vssd1 vssd1 vccd1 vccd1 _16798_/X sky130_fd_sc_hd__mux2_1
XFILLER_52_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18537_ _18542_/CLK _18537_/D vssd1 vssd1 vccd1 vccd1 _18537_/Q sky130_fd_sc_hd__dfxtp_2
X_15749_ _15754_/B _15746_/X _15748_/X _15740_/X vssd1 vssd1 vccd1 vccd1 _18516_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_209_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09270_ _09270_/A _09270_/B _09270_/C _09270_/D vssd1 vssd1 vccd1 vccd1 _09271_/C
+ sky130_fd_sc_hd__and4_1
X_18468_ _18469_/CLK _18468_/D vssd1 vssd1 vccd1 vccd1 _18468_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_205_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17419_ _17456_/A _17419_/B vssd1 vssd1 vccd1 vccd1 _17419_/Y sky130_fd_sc_hd__nand2_1
XFILLER_18_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18399_ _18404_/CLK _18399_/D vssd1 vssd1 vccd1 vccd1 _18399_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_193_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_193_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_228_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_228_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_195_wb_clk_i _18114_/CLK vssd1 vssd1 vccd1 vccd1 _18997_/CLK sky130_fd_sc_hd__clkbuf_16
Xclkbuf_leaf_124_wb_clk_i clkbuf_5_31_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18423_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_115_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_170_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_216_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08985_ _08985_/A vssd1 vssd1 vccd1 vccd1 _08985_/Y sky130_fd_sc_hd__inv_2
XFILLER_103_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_228_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19051__22 vssd1 vssd1 vccd1 vccd1 _19051__22/HI _19145_/A sky130_fd_sc_hd__conb_1
X_09606_ _10123_/A _10675_/A _09580_/A vssd1 vssd1 vccd1 vccd1 _09606_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_71_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_186_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_225_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09537_ _09568_/A _09537_/B vssd1 vssd1 vccd1 vccd1 _09540_/B sky130_fd_sc_hd__xor2_4
XFILLER_25_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_196_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09468_ _09468_/A vssd1 vssd1 vccd1 vccd1 _18136_/D sky130_fd_sc_hd__clkbuf_1
XPHY_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09399_ _18356_/Q _18355_/Q _18354_/Q vssd1 vssd1 vccd1 vccd1 _09402_/B sky130_fd_sc_hd__or3_4
XFILLER_138_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_1331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11430_ _17883_/Q vssd1 vssd1 vccd1 vccd1 _11431_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_71_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_138_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11361_ _11503_/A _11586_/C vssd1 vssd1 vccd1 vccd1 _11447_/A sky130_fd_sc_hd__nor2_1
XFILLER_137_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_125_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10312_ _10312_/A _10312_/B _10312_/C _09981_/A vssd1 vssd1 vccd1 vccd1 _10312_/X
+ sky130_fd_sc_hd__or4b_2
X_13100_ _13100_/A vssd1 vssd1 vccd1 vccd1 _18010_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_153_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14080_ _18734_/Q _13612_/X _13576_/X _18725_/Q _14079_/X vssd1 vssd1 vccd1 vccd1
+ _14080_/X sky130_fd_sc_hd__a221o_2
X_11292_ _11590_/B _11297_/C vssd1 vssd1 vccd1 vccd1 _11337_/A sky130_fd_sc_hd__nand2_1
XFILLER_106_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10243_ _10559_/S vssd1 vssd1 vccd1 vccd1 _10412_/A sky130_fd_sc_hd__buf_4
X_13031_ _17988_/Q _13015_/X _13030_/X vssd1 vssd1 vccd1 vccd1 _17988_/D sky130_fd_sc_hd__a21o_1
XFILLER_106_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10174_ _10547_/A vssd1 vssd1 vccd1 vccd1 _10939_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_152_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17770_ _19028_/Q _11040_/X _11035_/B _13381_/X _13339_/X vssd1 vssd1 vccd1 vccd1
+ _19028_/D sky130_fd_sc_hd__o2111a_1
X_14982_ _18371_/Q _18335_/Q _14994_/S vssd1 vssd1 vccd1 vccd1 _14982_/X sky130_fd_sc_hd__mux2_1
XFILLER_120_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16721_ _16723_/B _16719_/X _16720_/Y _16704_/X vssd1 vssd1 vccd1 vccd1 _18748_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_19_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13933_ _18319_/Q _13715_/X _13869_/A _18307_/Q _13932_/X vssd1 vssd1 vccd1 vccd1
+ _13933_/X sky130_fd_sc_hd__a221o_1
XFILLER_59_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16652_ _16678_/A _16796_/B _16652_/C vssd1 vssd1 vccd1 vccd1 _16652_/X sky130_fd_sc_hd__or3_1
X_13864_ _18838_/Q _13551_/X _13862_/X _13863_/X vssd1 vssd1 vccd1 vccd1 _13864_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_90_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_223_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15603_ _15605_/B _15601_/X _15602_/Y _15595_/X vssd1 vssd1 vccd1 vccd1 _18481_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_90_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12815_ _17960_/Q vssd1 vssd1 vccd1 vccd1 _12815_/Y sky130_fd_sc_hd__inv_2
XFILLER_216_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16583_ _17222_/A vssd1 vssd1 vccd1 vccd1 _16828_/A sky130_fd_sc_hd__clkbuf_2
X_13795_ _18297_/Q _13663_/X _13793_/X _13794_/X vssd1 vssd1 vccd1 vccd1 _13795_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_215_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18322_ _18350_/CLK _18322_/D vssd1 vssd1 vccd1 vccd1 _18322_/Q sky130_fd_sc_hd__dfxtp_4
X_15534_ _15570_/A _15534_/B vssd1 vssd1 vccd1 vccd1 _15534_/Y sky130_fd_sc_hd__nand2_1
XFILLER_203_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12746_ _12760_/A _12748_/A vssd1 vssd1 vccd1 vccd1 _12747_/B sky130_fd_sc_hd__nor2_1
XFILLER_43_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_203_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18253_ _18253_/CLK _18253_/D vssd1 vssd1 vccd1 vccd1 _18253_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15465_ _15529_/A vssd1 vssd1 vccd1 vccd1 _15599_/C sky130_fd_sc_hd__buf_2
XFILLER_175_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12677_ _17935_/Q vssd1 vssd1 vccd1 vccd1 _12691_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_30_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17204_ _18900_/Q _18864_/Q _17221_/S vssd1 vssd1 vccd1 vccd1 _17204_/X sky130_fd_sc_hd__mux2_1
XFILLER_187_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14416_ _09497_/B _14401_/X _14415_/Y vssd1 vssd1 vccd1 vccd1 _14417_/B sky130_fd_sc_hd__o21a_1
XFILLER_198_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11628_ _11614_/A _11615_/Y _11603_/B vssd1 vssd1 vccd1 vccd1 _11628_/Y sky130_fd_sc_hd__a21oi_1
X_18184_ _18184_/CLK _18184_/D vssd1 vssd1 vccd1 vccd1 _18184_/Q sky130_fd_sc_hd__dfxtp_2
X_15396_ _16909_/A vssd1 vssd1 vccd1 vccd1 _15997_/B sky130_fd_sc_hd__buf_2
XFILLER_128_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_204_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17135_ _18882_/Q _18846_/Q _17151_/S vssd1 vssd1 vccd1 vccd1 _17135_/X sky130_fd_sc_hd__mux2_1
XFILLER_50_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14347_ _14275_/A _14344_/X _14346_/X _14340_/X vssd1 vssd1 vccd1 vccd1 _18180_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_128_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11559_ _12267_/A _12261_/A _11645_/A _11556_/X _12274_/A vssd1 vssd1 vccd1 vccd1
+ _11559_/X sky130_fd_sc_hd__o311a_1
XFILLER_200_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17066_ _17068_/B _17064_/X _17065_/Y _17057_/X vssd1 vssd1 vccd1 vccd1 _18829_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_170_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14278_ _14319_/S _09915_/A _14277_/Y vssd1 vssd1 vccd1 vccd1 _14293_/A sky130_fd_sc_hd__a21oi_2
XFILLER_109_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16017_ _16064_/A _16017_/B vssd1 vssd1 vccd1 vccd1 _16017_/Y sky130_fd_sc_hd__nand2_1
X_13229_ _13233_/A _18070_/Q vssd1 vssd1 vccd1 vccd1 _13230_/A sky130_fd_sc_hd__and2_1
XFILLER_100_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_214_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17968_ _17969_/CLK _17968_/D vssd1 vssd1 vccd1 vccd1 _17968_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_66_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_226_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_214_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16919_ _16919_/A vssd1 vssd1 vccd1 vccd1 _17503_/A sky130_fd_sc_hd__buf_4
XFILLER_211_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17899_ _17901_/CLK _17899_/D vssd1 vssd1 vccd1 vccd1 _17899_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_66_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_211_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_226_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09322_ _09294_/X _09299_/X _09304_/X _09321_/Y vssd1 vssd1 vccd1 vccd1 _09339_/A
+ sky130_fd_sc_hd__a31o_1
XFILLER_55_1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_221_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09253_ _09253_/A _09253_/B _09253_/C _09253_/D vssd1 vssd1 vccd1 vccd1 _09254_/C
+ sky130_fd_sc_hd__and4_1
XFILLER_107_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_222_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09184_ _18602_/Q _18601_/Q _18600_/Q vssd1 vssd1 vccd1 vccd1 _09186_/C sky130_fd_sc_hd__or3_4
XFILLER_194_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_222_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_175_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08968_ _08972_/A vssd1 vssd1 vccd1 vccd1 _08968_/Y sky130_fd_sc_hd__inv_2
XTAP_4715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_229_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_216_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10930_ _10926_/X _10929_/X _10936_/S vssd1 vssd1 vccd1 vccd1 _10930_/X sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_92_wb_clk_i _18254_/CLK vssd1 vssd1 vccd1 vccd1 _18253_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_57_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_189_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_216_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10861_ _10833_/B _10853_/X _10860_/X vssd1 vssd1 vccd1 vccd1 _10861_/X sky130_fd_sc_hd__a21o_1
Xclkbuf_leaf_21_wb_clk_i clkbuf_5_4_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18902_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_186_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_231_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12600_ _12600_/A _12600_/B _12600_/C vssd1 vssd1 vccd1 vccd1 _12600_/Y sky130_fd_sc_hd__nand3_1
XPHY_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13580_ _13580_/A vssd1 vssd1 vccd1 vccd1 _13702_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_25_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10792_ _10838_/B _10778_/X _10787_/X _10791_/X _10622_/Y vssd1 vssd1 vccd1 vccd1
+ _10822_/A sky130_fd_sc_hd__o311a_1
XFILLER_231_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12531_ _12809_/A _12529_/X _12530_/Y vssd1 vssd1 vccd1 vccd1 _12531_/X sky130_fd_sc_hd__a21o_1
XFILLER_73_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_212_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15250_ _15250_/A vssd1 vssd1 vccd1 vccd1 _15267_/S sky130_fd_sc_hd__clkbuf_2
XPHY_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12462_ _12486_/B vssd1 vssd1 vccd1 vccd1 _12487_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_8_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14201_ _14297_/A _14355_/C _14355_/D _14463_/A vssd1 vssd1 vccd1 vccd1 _14275_/A
+ sky130_fd_sc_hd__o31a_1
XFILLER_71_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11413_ _11413_/A _11652_/A _11526_/B vssd1 vssd1 vccd1 vccd1 _11413_/Y sky130_fd_sc_hd__nor3b_2
X_15181_ _18419_/Q _18383_/Q _15198_/S vssd1 vssd1 vccd1 vccd1 _15181_/X sky130_fd_sc_hd__mux2_1
XFILLER_137_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12393_ _12394_/B _12394_/C _17896_/Q vssd1 vssd1 vccd1 vccd1 _12406_/A sky130_fd_sc_hd__o21a_1
XFILLER_201_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14132_ _18272_/Q _13507_/A _13500_/A _18296_/Q vssd1 vssd1 vccd1 vccd1 _14132_/X
+ sky130_fd_sc_hd__a22o_1
X_11344_ _17877_/Q _19030_/Q vssd1 vssd1 vccd1 vccd1 _11385_/A sky130_fd_sc_hd__or2b_1
XFILLER_152_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_1208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14063_ _18383_/Q _13546_/A _14059_/X _14062_/X vssd1 vssd1 vccd1 vccd1 _14063_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_153_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18940_ _18965_/CLK _18940_/D vssd1 vssd1 vccd1 vccd1 _18940_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_98_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11275_ _11806_/B _13442_/A vssd1 vssd1 vccd1 vccd1 _11275_/X sky130_fd_sc_hd__and2b_1
XFILLER_180_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13014_ _13041_/B vssd1 vssd1 vccd1 vccd1 _13025_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_80_1307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10226_ _10899_/A vssd1 vssd1 vccd1 vccd1 _11924_/A sky130_fd_sc_hd__buf_2
X_18871_ _18871_/CLK _18871_/D vssd1 vssd1 vccd1 vccd1 _18871_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_79_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17822_ _17824_/CLK _17822_/D vssd1 vssd1 vccd1 vccd1 _17822_/Q sky130_fd_sc_hd__dfxtp_1
X_10157_ _13389_/A _10137_/B _10135_/X vssd1 vssd1 vccd1 vccd1 _10165_/S sky130_fd_sc_hd__a21oi_2
XFILLER_94_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold4 hold4/A vssd1 vssd1 vccd1 vccd1 hold4/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_58_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14965_ _14975_/A _15257_/B _14965_/C vssd1 vssd1 vccd1 vccd1 _14965_/X sky130_fd_sc_hd__or3_1
X_17753_ _17753_/A vssd1 vssd1 vccd1 vccd1 _19019_/D sky130_fd_sc_hd__clkbuf_1
X_10088_ _09253_/C _09243_/C _10089_/S vssd1 vssd1 vccd1 vccd1 _10088_/X sky130_fd_sc_hd__mux2_1
XTAP_5994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13916_ _18769_/Q _14014_/A _14026_/A _18760_/Q vssd1 vssd1 vccd1 vccd1 _13916_/X
+ sky130_fd_sc_hd__a22o_1
X_16704_ _16760_/A vssd1 vssd1 vccd1 vccd1 _16704_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_48_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17684_ _17645_/X _17674_/Y _17675_/X _17676_/Y _18983_/Q vssd1 vssd1 vccd1 vccd1
+ _17685_/B sky130_fd_sc_hd__a32o_1
XFILLER_81_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_5_5_0_wb_clk_i clkbuf_5_5_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_5_5_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_2
X_14896_ _18349_/Q _18313_/Q _14905_/S vssd1 vssd1 vccd1 vccd1 _14896_/X sky130_fd_sc_hd__mux2_1
XFILLER_78_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16635_ _16634_/B _16633_/X _16634_/Y _16619_/X vssd1 vssd1 vccd1 vccd1 _18728_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_62_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13847_ _13847_/A vssd1 vssd1 vccd1 vccd1 _13848_/A sky130_fd_sc_hd__buf_8
XFILLER_74_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_223_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_204_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16566_ _16566_/A vssd1 vssd1 vccd1 vccd1 _16808_/A sky130_fd_sc_hd__buf_2
X_13778_ _18633_/Q _13749_/X _13774_/X _13777_/X vssd1 vssd1 vccd1 vccd1 _13778_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_62_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15517_ _15525_/B _15514_/X _15515_/X _15516_/X vssd1 vssd1 vccd1 vccd1 _18459_/D
+ sky130_fd_sc_hd__o211a_1
X_18305_ _18307_/CLK _18305_/D vssd1 vssd1 vccd1 vccd1 _18305_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_203_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12729_ _18095_/Q _12729_/B vssd1 vssd1 vccd1 vccd1 _12921_/A sky130_fd_sc_hd__nor2_1
XFILLER_31_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16497_ _16499_/B _16494_/X _16495_/Y _16496_/X vssd1 vssd1 vccd1 vccd1 _18694_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_148_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18236_ _18263_/CLK _18236_/D vssd1 vssd1 vccd1 vccd1 _18236_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15448_ _16041_/A _15448_/B vssd1 vssd1 vccd1 vccd1 _15460_/B sky130_fd_sc_hd__nor2_2
XFILLER_175_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_175_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_1272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18167_ _18967_/CLK _18167_/D vssd1 vssd1 vccd1 vccd1 _18167_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_102_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15379_ _18465_/Q _18429_/Q _15388_/S vssd1 vssd1 vccd1 vccd1 _15379_/X sky130_fd_sc_hd__mux2_1
XFILLER_144_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17118_ _17115_/B _17114_/X _17115_/Y _17117_/X vssd1 vssd1 vccd1 vccd1 _18842_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_85_1207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18098_ _18110_/CLK _18098_/D vssd1 vssd1 vccd1 vccd1 _18098_/Q sky130_fd_sc_hd__dfxtp_1
X_09940_ _10598_/A vssd1 vssd1 vccd1 vccd1 _10305_/S sky130_fd_sc_hd__buf_2
X_17049_ _18861_/Q _18825_/Q _17055_/S vssd1 vssd1 vccd1 vccd1 _17049_/X sky130_fd_sc_hd__mux2_1
XFILLER_217_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09871_ _09872_/A _09872_/B vssd1 vssd1 vccd1 vccd1 _09876_/B sky130_fd_sc_hd__xnor2_1
XTAP_731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_17 _09209_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_28 _09462_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_39 _10598_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_227_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_100_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_214_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_213_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_213_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09305_ _18455_/Q _18454_/Q _18453_/Q vssd1 vssd1 vccd1 vccd1 _09309_/A sky130_fd_sc_hd__or3_4
XFILLER_94_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_224_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_210_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09236_ _18944_/Q _18943_/Q _18942_/Q vssd1 vssd1 vccd1 vccd1 _09237_/D sky130_fd_sc_hd__or3_2
XFILLER_155_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_194_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_222_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09167_ _18650_/Q _18649_/Q _18648_/Q vssd1 vssd1 vccd1 vccd1 _09170_/B sky130_fd_sc_hd__or3_4
XFILLER_163_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09098_ _09098_/A _09098_/B _09098_/C _09098_/D vssd1 vssd1 vccd1 vccd1 _09104_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_107_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11060_ _17787_/Q vssd1 vssd1 vccd1 vccd1 _11336_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_153_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10011_ _09694_/A _10002_/X _10006_/X _10010_/X vssd1 vssd1 vccd1 vccd1 _10011_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_1_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_231_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14750_ _14750_/A _14753_/B vssd1 vssd1 vccd1 vccd1 _14750_/Y sky130_fd_sc_hd__nand2_1
XFILLER_218_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11962_ _12026_/B vssd1 vssd1 vccd1 vccd1 _12007_/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_3855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_229_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13701_ _18756_/Q _13856_/A _13493_/A _18747_/Q _13700_/X vssd1 vssd1 vccd1 vccd1
+ _13701_/X sky130_fd_sc_hd__a221o_1
XTAP_3866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_217_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10913_ _09319_/A _09309_/C _09314_/B _09319_/C _10430_/X _12032_/A vssd1 vssd1 vccd1
+ vccd1 _10914_/B sky130_fd_sc_hd__mux4_2
XTAP_3877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_205_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14681_ _14681_/A _14683_/B vssd1 vssd1 vccd1 vccd1 _14681_/Y sky130_fd_sc_hd__nand2_1
XTAP_3888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11893_ _17824_/Q _11891_/X _11892_/X vssd1 vssd1 vccd1 vccd1 _11893_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_72_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_229_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16420_ _16714_/A _16452_/B vssd1 vssd1 vccd1 vccd1 _16429_/B sky130_fd_sc_hd__nor2_1
X_13632_ _18462_/Q _13581_/X _13629_/X _13631_/X vssd1 vssd1 vccd1 vccd1 _13632_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_44_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10844_ _10700_/S _10838_/B _10842_/X _10843_/X vssd1 vssd1 vccd1 vccd1 _10844_/X
+ sky130_fd_sc_hd__o31a_1
XFILLER_220_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16351_ _16353_/B _16349_/X _16350_/Y _16334_/X vssd1 vssd1 vccd1 vccd1 _18658_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_164_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13563_ _13563_/A _13563_/B vssd1 vssd1 vccd1 vccd1 _13772_/A sky130_fd_sc_hd__nor2_1
X_10775_ _09304_/A _09294_/B _09299_/C _09304_/C _10687_/A _10770_/X vssd1 vssd1 vccd1
+ vccd1 _10775_/X sky130_fd_sc_hd__mux4_2
XFILLER_34_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_227_wb_clk_i _17864_/CLK vssd1 vssd1 vccd1 vccd1 _19035_/CLK sky130_fd_sc_hd__clkbuf_16
X_15302_ _18412_/Q _15303_/B _15301_/Y _15283_/X vssd1 vssd1 vccd1 vccd1 _18412_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_185_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12514_ _12514_/A vssd1 vssd1 vccd1 vccd1 _12514_/Y sky130_fd_sc_hd__inv_2
X_16282_ _18677_/Q _18641_/Q _16304_/S vssd1 vssd1 vccd1 vccd1 _16282_/X sky130_fd_sc_hd__mux2_1
XFILLER_160_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13494_ _13509_/B _13494_/B vssd1 vssd1 vccd1 vccd1 _13557_/A sky130_fd_sc_hd__nand2b_4
XFILLER_157_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18021_ _18095_/CLK _18021_/D vssd1 vssd1 vccd1 vccd1 _18021_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_8_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_199_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15233_ _15279_/A _15233_/B _15257_/C vssd1 vssd1 vccd1 vccd1 _15233_/X sky130_fd_sc_hd__or3_1
XFILLER_9_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12445_ _12437_/A _12438_/Y _12444_/Y vssd1 vssd1 vccd1 vccd1 _12452_/B sky130_fd_sc_hd__o21ai_1
X_15164_ _18415_/Q _18379_/Q _15177_/S vssd1 vssd1 vccd1 vccd1 _15164_/X sky130_fd_sc_hd__mux2_1
XFILLER_176_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12376_ _12365_/X _12369_/B _12375_/Y vssd1 vssd1 vccd1 vccd1 _12388_/B sky130_fd_sc_hd__a21oi_1
XFILLER_125_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14115_ _18932_/Q _13834_/X _13493_/X _18929_/Q _14114_/X vssd1 vssd1 vccd1 vccd1
+ _14115_/X sky130_fd_sc_hd__a221o_1
XFILLER_181_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11327_ _17876_/Q _17875_/Q vssd1 vssd1 vccd1 vccd1 _11339_/D sky130_fd_sc_hd__and2_1
XFILLER_99_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15095_ _15094_/B _15093_/X _15094_/Y _15083_/X vssd1 vssd1 vccd1 vccd1 _18362_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_141_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14046_ _18545_/Q _13697_/A _13537_/A _18521_/Q vssd1 vssd1 vccd1 vccd1 _14046_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_140_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18923_ _18959_/CLK _18923_/D vssd1 vssd1 vccd1 vccd1 _18923_/Q sky130_fd_sc_hd__dfxtp_4
X_11258_ _11501_/A _11258_/B _11584_/B vssd1 vssd1 vccd1 vccd1 _11586_/D sky130_fd_sc_hd__or3b_1
XFILLER_84_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10209_ _10210_/A _10210_/B vssd1 vssd1 vccd1 vccd1 _10211_/A sky130_fd_sc_hd__nor2_1
XFILLER_39_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18854_ _18862_/CLK _18854_/D vssd1 vssd1 vccd1 vccd1 _18854_/Q sky130_fd_sc_hd__dfxtp_4
X_11189_ _11190_/A _11196_/D vssd1 vssd1 vccd1 vccd1 _11191_/B sky130_fd_sc_hd__or2_1
XFILLER_68_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_227_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_209_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17805_ _17806_/CLK _17805_/D vssd1 vssd1 vccd1 vccd1 _17805_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15997_ _16043_/A _15997_/B _16021_/C vssd1 vssd1 vccd1 vccd1 _15997_/X sky130_fd_sc_hd__or3_1
X_18785_ _18785_/CLK _18785_/D vssd1 vssd1 vccd1 vccd1 _18785_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_5780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14948_ _14948_/A vssd1 vssd1 vccd1 vccd1 _14995_/A sky130_fd_sc_hd__buf_2
X_17736_ _17736_/A vssd1 vssd1 vccd1 vccd1 _17745_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_224_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XINSDIODE2_110 _14030_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14879_ _18345_/Q _18309_/Q _14883_/S vssd1 vssd1 vccd1 vccd1 _14879_/X sky130_fd_sc_hd__mux2_1
XFILLER_63_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17667_ _17667_/A vssd1 vssd1 vccd1 vccd1 _18978_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_208_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINSDIODE2_121 _15233_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XINSDIODE2_132 _15270_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_143 _17265_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16618_ _16631_/A _16623_/B vssd1 vssd1 vccd1 vccd1 _16618_/Y sky130_fd_sc_hd__nand2_1
XFILLER_211_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XINSDIODE2_154 _18387_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17598_ _17598_/A vssd1 vssd1 vccd1 vccd1 _18961_/D sky130_fd_sc_hd__clkbuf_1
XINSDIODE2_165 _18363_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_176 _18671_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16549_ _16621_/A vssd1 vssd1 vccd1 vccd1 _16565_/S sky130_fd_sc_hd__clkbuf_2
XINSDIODE2_187 _09103_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_198 _10434_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_210_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09021_ _09022_/A vssd1 vssd1 vccd1 vccd1 _09021_/Y sky130_fd_sc_hd__inv_2
XFILLER_136_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18219_ _18222_/CLK _18219_/D vssd1 vssd1 vccd1 vccd1 _18219_/Q sky130_fd_sc_hd__dfxtp_1
X_19199_ _19199_/A _08984_/Y vssd1 vssd1 vccd1 vccd1 io_out[37] sky130_fd_sc_hd__ebufn_8
XFILLER_129_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_191_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09923_ _09937_/A vssd1 vssd1 vccd1 vccd1 _09923_/X sky130_fd_sc_hd__buf_6
XFILLER_217_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09854_ _09866_/A _09866_/B _09853_/Y vssd1 vssd1 vccd1 vccd1 _09858_/B sky130_fd_sc_hd__o21ba_2
XFILLER_112_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_213_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_219_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09785_ _09792_/A _09785_/B vssd1 vssd1 vccd1 vccd1 _09785_/X sky130_fd_sc_hd__or2_1
XFILLER_100_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_214_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_230_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10560_ _09186_/C _09176_/B _10560_/S vssd1 vssd1 vccd1 vccd1 _10560_/X sky130_fd_sc_hd__mux2_1
XFILLER_10_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09219_ _09219_/A _09219_/B _09219_/C _09219_/D vssd1 vssd1 vccd1 vccd1 _09220_/C
+ sky130_fd_sc_hd__and4_1
X_10491_ _10484_/X _10491_/B vssd1 vssd1 vccd1 vccd1 _10491_/X sky130_fd_sc_hd__and2b_1
XFILLER_154_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12230_ _12517_/A _12230_/B vssd1 vssd1 vccd1 vccd1 _12231_/A sky130_fd_sc_hd__and2_1
XFILLER_68_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_182_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12161_ _17843_/Q _12172_/B vssd1 vssd1 vccd1 vccd1 _12161_/X sky130_fd_sc_hd__and2_1
XFILLER_146_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11112_ _11654_/B vssd1 vssd1 vccd1 vccd1 _13447_/A sky130_fd_sc_hd__buf_2
XFILLER_150_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12092_ _12092_/A _12092_/B vssd1 vssd1 vccd1 vccd1 _12092_/Y sky130_fd_sc_hd__nand2_1
XFILLER_151_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15920_ _18594_/Q _18558_/Q _15937_/S vssd1 vssd1 vccd1 vccd1 _15920_/X sky130_fd_sc_hd__mux2_1
XTAP_5010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11043_ _13368_/B vssd1 vssd1 vccd1 vccd1 _11044_/B sky130_fd_sc_hd__buf_2
XTAP_5021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_209_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15851_ _15853_/B _15849_/X _15850_/Y _15842_/X vssd1 vssd1 vccd1 vccd1 _18541_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_5054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14802_ _14814_/A _14802_/B vssd1 vssd1 vccd1 vccd1 _14802_/Y sky130_fd_sc_hd__nand2_1
XTAP_4364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15782_ _15818_/A _15782_/B vssd1 vssd1 vccd1 vccd1 _15782_/Y sky130_fd_sc_hd__nand2_1
X_18570_ _18577_/CLK _18570_/D vssd1 vssd1 vccd1 vccd1 _18570_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_40_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_224_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12994_ _10619_/A _12990_/A _12775_/A _12931_/A _17989_/Q vssd1 vssd1 vccd1 vccd1
+ _12994_/X sky130_fd_sc_hd__a32o_1
XFILLER_45_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14733_ _18309_/Q _18273_/Q _14736_/S vssd1 vssd1 vccd1 vccd1 _14733_/X sky130_fd_sc_hd__mux2_1
XFILLER_18_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17521_ _17541_/A _17524_/B vssd1 vssd1 vccd1 vccd1 _17521_/Y sky130_fd_sc_hd__nand2_1
XFILLER_205_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11945_ _11945_/A _11945_/B vssd1 vssd1 vccd1 vccd1 _11964_/C sky130_fd_sc_hd__nand2_1
XFILLER_44_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17452_ _18961_/Q _18925_/Q _17467_/S vssd1 vssd1 vccd1 vccd1 _17452_/X sky130_fd_sc_hd__mux2_1
XTAP_2962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14664_ _16935_/A vssd1 vssd1 vccd1 vccd1 _15257_/B sky130_fd_sc_hd__buf_6
XFILLER_178_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11876_ _18164_/Q _11867_/X _11875_/Y vssd1 vssd1 vccd1 vccd1 _11877_/B sky130_fd_sc_hd__a21oi_1
XTAP_2984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_229_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16403_ _16407_/B _16400_/X _16402_/Y _16398_/X vssd1 vssd1 vccd1 vccd1 _18670_/D
+ sky130_fd_sc_hd__o211a_1
X_13615_ _13615_/A vssd1 vssd1 vccd1 vccd1 _13616_/A sky130_fd_sc_hd__buf_6
XFILLER_220_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17383_ _17395_/A _17383_/B vssd1 vssd1 vccd1 vccd1 _17383_/Y sky130_fd_sc_hd__nand2_1
X_10827_ _09227_/D _10644_/A _10826_/X _10852_/A vssd1 vssd1 vccd1 vccd1 _10827_/X
+ sky130_fd_sc_hd__o211a_1
X_14595_ _14651_/A _15197_/A vssd1 vssd1 vccd1 vccd1 _14606_/B sky130_fd_sc_hd__nor2_2
XFILLER_125_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16334_ _16354_/A vssd1 vssd1 vccd1 vccd1 _16334_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_199_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13546_ _13546_/A vssd1 vssd1 vccd1 vccd1 _13546_/X sky130_fd_sc_hd__clkbuf_4
X_10758_ _09309_/A _10575_/A _09319_/D _09309_/D _10693_/X _10660_/X vssd1 vssd1 vccd1
+ vccd1 _10758_/X sky130_fd_sc_hd__mux4_1
XFILLER_185_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16265_ _16265_/A _16268_/B vssd1 vssd1 vccd1 vccd1 _16265_/Y sky130_fd_sc_hd__nand2_1
XFILLER_187_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13477_ _17846_/Q _13457_/X _13465_/X vssd1 vssd1 vccd1 vccd1 _13478_/B sky130_fd_sc_hd__a21oi_1
X_10689_ _10689_/A _10838_/B _10689_/C vssd1 vssd1 vccd1 vccd1 _10689_/X sky130_fd_sc_hd__and3_1
X_15216_ _15239_/A _15216_/B vssd1 vssd1 vccd1 vccd1 _15216_/Y sky130_fd_sc_hd__nand2_1
X_18004_ _18997_/CLK _18004_/D vssd1 vssd1 vccd1 vccd1 _18004_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_195_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_145_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12428_ _12426_/B _12426_/C _17900_/Q vssd1 vssd1 vccd1 vccd1 _12439_/B sky130_fd_sc_hd__a21bo_1
X_16196_ _16202_/B _16192_/X _16195_/X _16185_/X vssd1 vssd1 vccd1 vccd1 _18621_/D
+ sky130_fd_sc_hd__o211a_1
X_15147_ _15292_/A _15279_/C vssd1 vssd1 vccd1 vccd1 _15154_/B sky130_fd_sc_hd__nor2_2
XFILLER_142_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12359_ _12352_/B _12493_/B _14457_/B _17892_/Q vssd1 vssd1 vccd1 vccd1 _12359_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_153_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15078_ _18394_/Q _18358_/Q _15081_/S vssd1 vssd1 vccd1 vccd1 _15078_/X sky130_fd_sc_hd__mux2_1
XFILLER_142_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14029_ _18254_/Q _13856_/X _13858_/X _18245_/Q _14028_/X vssd1 vssd1 vccd1 vccd1
+ _14029_/X sky130_fd_sc_hd__a221o_1
X_18906_ _18908_/CLK _18906_/D vssd1 vssd1 vccd1 vccd1 _18906_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_68_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18837_ _18875_/CLK _18837_/D vssd1 vssd1 vccd1 vccd1 _18837_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_222_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09570_ _10142_/A _09570_/B vssd1 vssd1 vccd1 vccd1 _09570_/X sky130_fd_sc_hd__or2_1
X_18768_ _18773_/CLK _18768_/D vssd1 vssd1 vccd1 vccd1 _18768_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_208_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_224_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17719_ _17723_/A _19005_/Q vssd1 vssd1 vccd1 vccd1 _17720_/A sky130_fd_sc_hd__and2_1
X_18699_ _18701_/CLK _18699_/D vssd1 vssd1 vccd1 vccd1 _18699_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_224_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_149_wb_clk_i clkbuf_5_26_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18307_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_63_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_196_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_220_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_1295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_177_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_178_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09004_ input1/X vssd1 vssd1 vccd1 vccd1 _09029_/A sky130_fd_sc_hd__buf_4
XFILLER_178_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_191_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_219_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_219_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09906_ _09365_/B _09370_/C _09365_/D _09360_/D _10274_/S _09905_/X vssd1 vssd1 vccd1
+ vccd1 _09906_/X sky130_fd_sc_hd__mux4_1
XFILLER_160_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_1282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09837_ _13348_/A _10629_/A vssd1 vssd1 vccd1 vccd1 _09837_/Y sky130_fd_sc_hd__nand2_1
XFILLER_219_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_189_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09768_ _18115_/Q vssd1 vssd1 vccd1 vccd1 _09781_/A sky130_fd_sc_hd__clkinv_2
XFILLER_206_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09699_ _12078_/A _09699_/B vssd1 vssd1 vccd1 vccd1 _10024_/A sky130_fd_sc_hd__xnor2_4
XTAP_2236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_199_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11730_ _11730_/A _11730_/B vssd1 vssd1 vccd1 vccd1 _11730_/Y sky130_fd_sc_hd__nand2_1
XTAP_1524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_214_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11661_ _11661_/A _11665_/B vssd1 vssd1 vccd1 vccd1 _11669_/B sky130_fd_sc_hd__or2_1
XFILLER_35_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13400_ _09822_/A _13368_/A _13368_/B _13386_/Y vssd1 vssd1 vccd1 vccd1 _13401_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_186_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10612_ _10612_/A _10612_/B _18121_/Q vssd1 vssd1 vccd1 vccd1 _10731_/B sky130_fd_sc_hd__nor3b_4
XFILLER_211_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14380_ _14373_/A _14373_/B _15015_/B vssd1 vssd1 vccd1 vccd1 _14381_/B sky130_fd_sc_hd__a21oi_1
X_11592_ _11899_/C _11808_/B _11592_/C _11592_/D vssd1 vssd1 vccd1 vccd1 _11868_/B
+ sky130_fd_sc_hd__nor4_4
XFILLER_10_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13331_ _18094_/Q _13329_/X _13330_/Y vssd1 vssd1 vccd1 vccd1 _18094_/D sky130_fd_sc_hd__o21ai_1
XFILLER_35_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10543_ _09386_/A _09376_/B _09381_/C _09972_/A _10518_/A _10542_/X vssd1 vssd1 vccd1
+ vccd1 _10543_/X sky130_fd_sc_hd__mux4_1
XFILLER_194_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_202_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16050_ _18626_/Q _18590_/Q _16050_/S vssd1 vssd1 vccd1 vccd1 _16050_/X sky130_fd_sc_hd__mux2_1
XFILLER_143_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13262_ _13266_/A _18085_/Q vssd1 vssd1 vccd1 vccd1 _13263_/A sky130_fd_sc_hd__and2_1
XFILLER_108_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10474_ _10902_/S _10474_/B vssd1 vssd1 vccd1 vccd1 _10474_/X sky130_fd_sc_hd__or2_1
XFILLER_183_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15001_ _15134_/B vssd1 vssd1 vccd1 vccd1 _15054_/C sky130_fd_sc_hd__clkbuf_2
X_12213_ _12257_/A vssd1 vssd1 vccd1 vccd1 _14504_/B sky130_fd_sc_hd__buf_8
XFILLER_170_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13193_ _13197_/A _18054_/Q vssd1 vssd1 vccd1 vccd1 _13194_/A sky130_fd_sc_hd__and2_1
XFILLER_135_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12144_ _17943_/Q _18167_/Q _12144_/S vssd1 vssd1 vccd1 vccd1 _12145_/A sky130_fd_sc_hd__mux2_2
XFILLER_124_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16952_ _16952_/A vssd1 vssd1 vccd1 vccd1 _16970_/S sky130_fd_sc_hd__clkbuf_2
X_12075_ _13372_/A _10829_/X _13353_/A vssd1 vssd1 vccd1 vccd1 _12075_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_1_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11026_ _11026_/A vssd1 vssd1 vccd1 vccd1 _11026_/X sky130_fd_sc_hd__buf_2
X_15903_ _17119_/A _17119_/B _15903_/C _16512_/C vssd1 vssd1 vccd1 vccd1 _16366_/B
+ sky130_fd_sc_hd__or4b_4
XFILLER_133_1355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16883_ _18787_/Q _16884_/B _16882_/Y _16871_/X vssd1 vssd1 vccd1 vccd1 _18787_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_38_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18622_ _18623_/CLK _18622_/D vssd1 vssd1 vccd1 vccd1 _18622_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_92_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15834_ _15839_/B _15832_/X _15833_/X _15823_/X vssd1 vssd1 vccd1 vccd1 _18537_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_4150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_225_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18553_ _18553_/CLK _18553_/D vssd1 vssd1 vccd1 vccd1 _18553_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15765_ _15885_/A vssd1 vssd1 vccd1 vccd1 _15815_/A sky130_fd_sc_hd__clkbuf_2
XTAP_3460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12977_ _12976_/A _12976_/B _12962_/A vssd1 vssd1 vccd1 vccd1 _12977_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_206_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17504_ _18975_/Q _18939_/Q _17515_/S vssd1 vssd1 vccd1 vccd1 _17504_/X sky130_fd_sc_hd__mux2_1
X_14716_ _14778_/A vssd1 vssd1 vccd1 vccd1 _14716_/X sky130_fd_sc_hd__clkbuf_2
X_11928_ _11932_/A _11930_/B _12021_/A vssd1 vssd1 vccd1 vccd1 _11945_/B sky130_fd_sc_hd__a21o_1
XFILLER_75_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18484_ _18485_/CLK _18484_/D vssd1 vssd1 vccd1 vccd1 _18484_/Q sky130_fd_sc_hd__dfxtp_2
X_15696_ _15993_/A _15696_/B vssd1 vssd1 vccd1 vccd1 _15708_/B sky130_fd_sc_hd__nor2_1
XTAP_2770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_177_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14647_ _14668_/A vssd1 vssd1 vccd1 vccd1 _14647_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_127_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17435_ _17435_/A _17491_/B vssd1 vssd1 vccd1 vccd1 _17444_/B sky130_fd_sc_hd__nor2_2
XFILLER_166_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11859_ _11859_/A vssd1 vssd1 vccd1 vccd1 _11860_/B sky130_fd_sc_hd__inv_2
XFILLER_53_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_220_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14578_ _14685_/B vssd1 vssd1 vccd1 vccd1 _17687_/B sky130_fd_sc_hd__buf_2
X_17366_ _17372_/B _17364_/X _17365_/X _17361_/X vssd1 vssd1 vccd1 vccd1 _18903_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_203_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_220_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16317_ _16329_/A _16317_/B vssd1 vssd1 vccd1 vccd1 _16317_/Y sky130_fd_sc_hd__nand2_1
X_13529_ _13529_/A vssd1 vssd1 vccd1 vccd1 _13731_/A sky130_fd_sc_hd__buf_4
XFILLER_174_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17297_ _17303_/B _17295_/X _17296_/X _17283_/X vssd1 vssd1 vccd1 vccd1 _18885_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_158_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19127__98 vssd1 vssd1 vccd1 vccd1 _19127__98/HI _19235_/A sky130_fd_sc_hd__conb_1
X_16248_ _16248_/A _16692_/B _16272_/C vssd1 vssd1 vccd1 vccd1 _16248_/X sky130_fd_sc_hd__or3_1
XFILLER_174_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16179_ _18654_/Q _18618_/Q _16192_/S vssd1 vssd1 vccd1 vccd1 _16179_/X sky130_fd_sc_hd__mux2_1
XFILLER_154_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_217_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_1305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_228_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09622_ _10204_/A _17975_/Q vssd1 vssd1 vccd1 vccd1 _09623_/B sky130_fd_sc_hd__xor2_2
XFILLER_216_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09553_ _10123_/A _10114_/B vssd1 vssd1 vccd1 vccd1 _09553_/Y sky130_fd_sc_hd__nand2_1
XFILLER_71_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09484_ _18146_/D _09463_/A _09461_/A _18150_/D vssd1 vssd1 vccd1 vccd1 _18149_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_23_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_224_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_212_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_211_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_212_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_177_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_221_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_178_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_46_wb_clk_i clkbuf_5_5_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18871_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_164_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_1333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10190_ _18120_/Q _10193_/B _09837_/Y vssd1 vssd1 vccd1 vccd1 _10258_/B sky130_fd_sc_hd__a21bo_1
XFILLER_219_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_1366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12900_ _17963_/Q _12899_/B _12854_/X vssd1 vssd1 vccd1 vccd1 _12901_/B sky130_fd_sc_hd__o21ai_1
XFILLER_87_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_219_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13880_ _18910_/Q _13657_/X _13731_/A _18904_/Q vssd1 vssd1 vccd1 vccd1 _13880_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_189_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_228_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12831_ _12646_/A _12792_/X _17965_/Q _12697_/B _12830_/X vssd1 vssd1 vccd1 vccd1
+ _12835_/C sky130_fd_sc_hd__a221o_1
XTAP_2011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15550_ _18504_/Q _18468_/Q _15565_/S vssd1 vssd1 vccd1 vccd1 _15550_/X sky130_fd_sc_hd__mux2_1
XTAP_2044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12762_ _18151_/Q _12721_/X _13271_/A _12761_/X vssd1 vssd1 vccd1 vccd1 _12762_/X
+ sky130_fd_sc_hd__o31a_1
XTAP_2055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14501_ _14501_/A vssd1 vssd1 vccd1 vccd1 _18224_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11713_ _11253_/A _11712_/X _11683_/C _11595_/Y vssd1 vssd1 vccd1 vccd1 _11714_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_14_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15481_ _15492_/A _15921_/B _15515_/C vssd1 vssd1 vccd1 vccd1 _15481_/X sky130_fd_sc_hd__or3_1
XTAP_2099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12693_ _12693_/A _12693_/B vssd1 vssd1 vccd1 vccd1 _12693_/Y sky130_fd_sc_hd__nand2_1
XTAP_1376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_202_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14432_ _18198_/Q _14431_/X _14428_/X _09501_/B vssd1 vssd1 vccd1 vccd1 _14433_/B
+ sky130_fd_sc_hd__o2bb2a_1
X_17220_ _17230_/B _17216_/X _17217_/X _17219_/X vssd1 vssd1 vccd1 vccd1 _18867_/D
+ sky130_fd_sc_hd__o211a_1
X_11644_ _17861_/Q _11671_/B vssd1 vssd1 vccd1 vccd1 _11673_/A sky130_fd_sc_hd__or2_1
XFILLER_230_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17151_ _18886_/Q _18850_/Q _17151_/S vssd1 vssd1 vccd1 vccd1 _17151_/X sky130_fd_sc_hd__mux2_1
X_14363_ _14422_/A _14510_/B _13416_/A vssd1 vssd1 vccd1 vccd1 _14373_/C sky130_fd_sc_hd__a21oi_1
X_11575_ _11553_/Y _11390_/A _11525_/B _11570_/B vssd1 vssd1 vccd1 vccd1 _11575_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_10_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16102_ _16853_/A vssd1 vssd1 vccd1 vccd1 _16703_/B sky130_fd_sc_hd__buf_4
XFILLER_156_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_196_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13314_ _13314_/A vssd1 vssd1 vccd1 vccd1 _13324_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_17082_ _17514_/A _17107_/B vssd1 vssd1 vccd1 vccd1 _17091_/B sky130_fd_sc_hd__nor2_2
X_10526_ _10520_/X _10525_/X _10936_/S vssd1 vssd1 vccd1 vccd1 _10526_/X sky130_fd_sc_hd__mux2_1
XFILLER_182_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14294_ _14311_/A _14294_/B vssd1 vssd1 vccd1 vccd1 _14294_/X sky130_fd_sc_hd__or2_1
XFILLER_7_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16033_ _16039_/B _16031_/X _16032_/X _16028_/X vssd1 vssd1 vccd1 vccd1 _18585_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_171_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_170_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13245_ _13245_/A vssd1 vssd1 vccd1 vccd1 _18076_/D sky130_fd_sc_hd__clkbuf_1
X_10457_ _10542_/A vssd1 vssd1 vccd1 vccd1 _10484_/A sky130_fd_sc_hd__buf_4
XFILLER_100_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13176_ _13176_/A vssd1 vssd1 vccd1 vccd1 _18045_/D sky130_fd_sc_hd__clkbuf_1
X_10388_ _10388_/A _10388_/B vssd1 vssd1 vccd1 vccd1 _10388_/X sky130_fd_sc_hd__or2_1
XFILLER_151_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12127_ _12127_/A _12127_/B _12127_/C _12127_/D vssd1 vssd1 vccd1 vccd1 _12132_/A
+ sky130_fd_sc_hd__or4_1
XFILLER_151_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17984_ _17987_/CLK _17984_/D vssd1 vssd1 vccd1 vccd1 _17984_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_123_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16935_ _16935_/A vssd1 vssd1 vccd1 vccd1 _17516_/B sky130_fd_sc_hd__buf_6
XFILLER_81_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12058_ _12059_/A _13526_/A vssd1 vssd1 vccd1 vccd1 _12058_/X sky130_fd_sc_hd__or2_1
XFILLER_77_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11009_ _17807_/Q vssd1 vssd1 vccd1 vccd1 _11181_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_133_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16866_ _16866_/A _17460_/B _16866_/C vssd1 vssd1 vccd1 vccd1 _16866_/X sky130_fd_sc_hd__or3_1
XFILLER_92_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18605_ _18607_/CLK _18605_/D vssd1 vssd1 vccd1 vccd1 _18605_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_19_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_225_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15817_ _18569_/Q _18533_/Q _15838_/S vssd1 vssd1 vccd1 vccd1 _15817_/X sky130_fd_sc_hd__mux2_1
XFILLER_203_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16797_ _16803_/B _16795_/X _16796_/X _16781_/X vssd1 vssd1 vccd1 vccd1 _18768_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_53_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18536_ _18546_/CLK _18536_/D vssd1 vssd1 vccd1 vccd1 _18536_/Q sky130_fd_sc_hd__dfxtp_1
X_15748_ _15799_/A _16043_/B _15748_/C vssd1 vssd1 vccd1 vccd1 _15748_/X sky130_fd_sc_hd__or3_1
XTAP_3290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_221_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18467_ _18467_/CLK _18467_/D vssd1 vssd1 vccd1 vccd1 _18467_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_61_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15679_ _18498_/Q _15683_/B _15678_/X _15662_/X vssd1 vssd1 vccd1 vccd1 _18498_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_209_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17418_ _18916_/Q _17419_/B _17417_/Y _17400_/X vssd1 vssd1 vccd1 vccd1 _18916_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_21_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_221_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18398_ _18398_/CLK _18398_/D vssd1 vssd1 vccd1 vccd1 _18398_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_194_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_187_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17349_ _17395_/A _17349_/B vssd1 vssd1 vccd1 vccd1 _17349_/Y sky130_fd_sc_hd__nand2_1
XFILLER_9_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_1355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_228_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19019_ _19019_/CLK _19019_/D vssd1 vssd1 vccd1 vccd1 _19019_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_115_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_216_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08984_ _08985_/A vssd1 vssd1 vccd1 vccd1 _08984_/Y sky130_fd_sc_hd__inv_2
XFILLER_87_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_1271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_164_wb_clk_i clkbuf_5_10_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18069_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_56_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09605_ _10155_/C vssd1 vssd1 vccd1 vccd1 _10675_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_113_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_228_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_227_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09536_ _09565_/A _10114_/B vssd1 vssd1 vccd1 vccd1 _09537_/B sky130_fd_sc_hd__xnor2_2
XFILLER_71_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_227_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_184_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09467_ _09467_/A _09467_/B vssd1 vssd1 vccd1 vccd1 _09468_/A sky130_fd_sc_hd__or2_1
XFILLER_58_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_196_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09398_ _18353_/Q _18352_/Q _18351_/Q vssd1 vssd1 vccd1 vccd1 _09402_/A sky130_fd_sc_hd__or3_2
XFILLER_11_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_138_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11360_ _11506_/B vssd1 vssd1 vccd1 vccd1 _11586_/C sky130_fd_sc_hd__clkinv_2
XFILLER_164_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10311_ _10305_/S _10306_/X _10310_/X _09930_/A vssd1 vssd1 vccd1 vccd1 _10312_/C
+ sky130_fd_sc_hd__o211a_1
XFILLER_4_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11291_ _17787_/Q _17786_/Q _17785_/Q _11334_/B vssd1 vssd1 vccd1 vccd1 _11297_/C
+ sky130_fd_sc_hd__a31o_1
XFILLER_180_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13030_ _13016_/X _12990_/A _12935_/X _13210_/A vssd1 vssd1 vccd1 vccd1 _13030_/X
+ sky130_fd_sc_hd__a31o_1
X_10242_ _10561_/S vssd1 vssd1 vccd1 vccd1 _10498_/A sky130_fd_sc_hd__buf_2
XFILLER_69_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10173_ _12053_/A _12053_/B vssd1 vssd1 vccd1 vccd1 _10547_/A sky130_fd_sc_hd__nand2_2
XFILLER_152_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14981_ _14983_/B _14978_/X _14979_/Y _14980_/X vssd1 vssd1 vccd1 vccd1 _18334_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_94_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_208_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16720_ _16752_/A _16723_/B vssd1 vssd1 vccd1 vccd1 _16720_/Y sky130_fd_sc_hd__nand2_1
X_13932_ _18313_/Q _13734_/A _13721_/X _18331_/Q vssd1 vssd1 vccd1 vccd1 _13932_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_120_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16651_ _18768_/Q _18732_/Q _16657_/S vssd1 vssd1 vccd1 vccd1 _16651_/X sky130_fd_sc_hd__mux2_1
X_13863_ _18826_/Q _13596_/X _13630_/X _18808_/Q vssd1 vssd1 vccd1 vccd1 _13863_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_130_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15602_ _15630_/A _15605_/B vssd1 vssd1 vccd1 vccd1 _15602_/Y sky130_fd_sc_hd__nand2_1
X_12814_ _12653_/B _17959_/Q _12794_/X _12797_/X _12813_/X vssd1 vssd1 vccd1 vccd1
+ _12814_/X sky130_fd_sc_hd__a2111o_1
XFILLER_222_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16582_ _18714_/Q _16589_/B _16579_/X _16581_/X vssd1 vssd1 vccd1 vccd1 _18714_/D
+ sky130_fd_sc_hd__o211a_1
X_13794_ _18285_/Q _13785_/X _13766_/X _18267_/Q vssd1 vssd1 vccd1 vccd1 _13794_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_188_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_216_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18321_ _18350_/CLK _18321_/D vssd1 vssd1 vccd1 vccd1 _18321_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_231_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15533_ _18463_/Q _15534_/B _15532_/Y _15516_/X vssd1 vssd1 vccd1 vccd1 _18463_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_1140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12745_ _18993_/Q vssd1 vssd1 vccd1 vccd1 _12760_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_203_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15464_ _15757_/A _17265_/A vssd1 vssd1 vccd1 vccd1 _15529_/A sky130_fd_sc_hd__or2_2
X_18252_ _18253_/CLK _18252_/D vssd1 vssd1 vccd1 vccd1 _18252_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12676_ _17936_/Q _12676_/B vssd1 vssd1 vccd1 vccd1 _12679_/A sky130_fd_sc_hd__xnor2_1
XFILLER_175_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14415_ _14405_/X _14414_/Y _18194_/Q vssd1 vssd1 vccd1 vccd1 _14415_/Y sky130_fd_sc_hd__o21ai_1
X_17203_ _17226_/A vssd1 vssd1 vccd1 vccd1 _17221_/S sky130_fd_sc_hd__clkbuf_2
X_11627_ _11615_/Y _11626_/X _11603_/Y vssd1 vssd1 vccd1 vccd1 _11627_/Y sky130_fd_sc_hd__a21boi_1
XFILLER_50_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15395_ _18468_/Q _18432_/Q _15412_/S vssd1 vssd1 vccd1 vccd1 _15395_/X sky130_fd_sc_hd__mux2_1
X_18183_ _18184_/CLK _18183_/D vssd1 vssd1 vccd1 vccd1 _18183_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_30_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14346_ _14299_/X _14272_/B _14283_/A _14300_/X _17119_/A vssd1 vssd1 vccd1 vccd1
+ _14346_/X sky130_fd_sc_hd__a311o_1
X_17134_ _17226_/A vssd1 vssd1 vccd1 vccd1 _17151_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_204_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11558_ _11562_/A _12269_/A vssd1 vssd1 vccd1 vccd1 _12274_/A sky130_fd_sc_hd__nand2_1
XFILLER_129_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_183_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10509_ _09153_/B _09993_/A _10509_/S vssd1 vssd1 vccd1 vccd1 _10509_/X sky130_fd_sc_hd__mux2_1
X_17065_ _17088_/A _17068_/B vssd1 vssd1 vccd1 vccd1 _17065_/Y sky130_fd_sc_hd__nand2_1
X_14277_ _12031_/A _14205_/A _14276_/X vssd1 vssd1 vccd1 vccd1 _14277_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_195_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11489_ _17888_/Q _11489_/B vssd1 vssd1 vccd1 vccd1 _12336_/B sky130_fd_sc_hd__and2_1
XFILLER_48_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16016_ _16216_/A vssd1 vssd1 vccd1 vccd1 _16064_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_170_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13228_ _13228_/A vssd1 vssd1 vccd1 vccd1 _18068_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_170_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13159_ _13159_/A vssd1 vssd1 vccd1 vccd1 _18037_/D sky130_fd_sc_hd__clkbuf_1
XTAP_924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17967_ _17969_/CLK _17967_/D vssd1 vssd1 vccd1 vccd1 _17967_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_97_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16918_ _16916_/B _16915_/X _16916_/Y _16917_/X vssd1 vssd1 vccd1 vccd1 _18794_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_226_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17898_ _17901_/CLK _17898_/D vssd1 vssd1 vccd1 vccd1 _17898_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_93_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_0_wb_clk_i wb_clk_i vssd1 vssd1 vccd1 vccd1 clkbuf_0_wb_clk_i/X sky130_fd_sc_hd__clkbuf_16
X_16849_ _16847_/B _16846_/X _16847_/Y _16848_/X vssd1 vssd1 vccd1 vccd1 _18779_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_93_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_214_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_226_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_225_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_213_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09321_ _09321_/A vssd1 vssd1 vccd1 vccd1 _09321_/Y sky130_fd_sc_hd__inv_2
XFILLER_34_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18519_ _18546_/CLK _18519_/D vssd1 vssd1 vccd1 vccd1 _18519_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_146_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09252_ _18911_/Q _18910_/Q _18909_/Q vssd1 vssd1 vccd1 vccd1 _09253_/D sky130_fd_sc_hd__or3_4
XFILLER_221_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_193_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_178_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09183_ _18623_/Q _18622_/Q _18621_/Q vssd1 vssd1 vccd1 vccd1 _09186_/B sky130_fd_sc_hd__or3_4
XFILLER_18_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_222_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_193_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_222_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_190_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19111__82 vssd1 vssd1 vccd1 vccd1 _19111__82/HI _19219_/A sky130_fd_sc_hd__conb_1
XTAP_5417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08967_ _08967_/A vssd1 vssd1 vccd1 vccd1 _08972_/A sky130_fd_sc_hd__buf_12
XTAP_5439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_229_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10860_ _10616_/Y _10856_/X _10859_/X _10733_/X vssd1 vssd1 vccd1 vccd1 _10860_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_72_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_216_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09519_ _17780_/Q _09509_/Y _09518_/X _17779_/Q vssd1 vssd1 vccd1 vccd1 _17779_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_231_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_140_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10791_ _10779_/X _10843_/C _10788_/X _10790_/X _10671_/B vssd1 vssd1 vccd1 vccd1
+ _10791_/X sky130_fd_sc_hd__a311o_1
XPHY_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_227_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12530_ _17916_/Q vssd1 vssd1 vccd1 vccd1 _12530_/Y sky130_fd_sc_hd__inv_2
XPHY_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_61_wb_clk_i _18759_/CLK vssd1 vssd1 vccd1 vccd1 _18722_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_169_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_185_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12461_ _12477_/A _12477_/B vssd1 vssd1 vccd1 vccd1 _12466_/B sky130_fd_sc_hd__or2_1
XFILLER_36_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14200_ _14300_/A vssd1 vssd1 vccd1 vccd1 _14463_/A sky130_fd_sc_hd__inv_2
X_11412_ _11412_/A _11732_/A _11412_/C _11594_/A vssd1 vssd1 vccd1 vccd1 _11526_/B
+ sky130_fd_sc_hd__or4_2
XFILLER_201_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15180_ _15250_/A vssd1 vssd1 vccd1 vccd1 _15198_/S sky130_fd_sc_hd__clkbuf_2
X_12392_ _12384_/B _18988_/Q vssd1 vssd1 vccd1 vccd1 _12394_/C sky130_fd_sc_hd__and2b_1
XFILLER_123_1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14131_ _18287_/Q _14124_/A _13706_/X _18269_/Q vssd1 vssd1 vccd1 vccd1 _14131_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_125_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11343_ _17878_/Q vssd1 vssd1 vccd1 vccd1 _11346_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_192_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14062_ _18407_/Q _13940_/X _14060_/X _14061_/X vssd1 vssd1 vccd1 vccd1 _14062_/X
+ sky130_fd_sc_hd__a211o_1
X_11274_ _17787_/Q _17786_/Q _17785_/Q vssd1 vssd1 vccd1 vccd1 _11806_/B sky130_fd_sc_hd__nor3_2
XFILLER_140_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13013_ _18151_/Q _13019_/B vssd1 vssd1 vccd1 vccd1 _13041_/B sky130_fd_sc_hd__nand2_1
X_10225_ _10555_/A vssd1 vssd1 vccd1 vccd1 _10899_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_79_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18870_ _18870_/CLK _18870_/D vssd1 vssd1 vccd1 vccd1 _18870_/Q sky130_fd_sc_hd__dfxtp_2
X_17821_ _17821_/CLK _17821_/D vssd1 vssd1 vccd1 vccd1 _17821_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_95_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10156_ _10169_/A _10154_/X _10155_/X vssd1 vssd1 vccd1 vccd1 _10158_/A sky130_fd_sc_hd__a21oi_1
XFILLER_94_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_181_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17752_ _17756_/A _19020_/Q vssd1 vssd1 vccd1 vccd1 _17753_/A sky130_fd_sc_hd__and2_1
XFILLER_48_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14964_ _18366_/Q _18330_/Q _14974_/S vssd1 vssd1 vccd1 vccd1 _14964_/X sky130_fd_sc_hd__mux2_1
XFILLER_134_1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10087_ _09270_/A _10813_/A _09265_/C _09265_/A _10102_/S _10090_/S vssd1 vssd1 vccd1
+ vccd1 _10087_/X sky130_fd_sc_hd__mux4_1
XTAP_5984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16703_ _16736_/A _16703_/B _16716_/C vssd1 vssd1 vccd1 vccd1 _16703_/X sky130_fd_sc_hd__or3_1
XFILLER_47_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13915_ _13649_/X _13890_/X _13914_/X _14507_/B vssd1 vssd1 vccd1 vccd1 _13915_/X
+ sky130_fd_sc_hd__a211o_1
X_17683_ _17736_/A vssd1 vssd1 vccd1 vccd1 _17712_/A sky130_fd_sc_hd__buf_4
X_14895_ _14900_/B _14893_/X _14894_/X _14881_/X vssd1 vssd1 vccd1 vccd1 _18312_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_48_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16634_ _16634_/A _16634_/B vssd1 vssd1 vccd1 vccd1 _16634_/Y sky130_fd_sc_hd__nand2_1
XFILLER_90_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13846_ _13836_/X _13845_/X _12042_/B vssd1 vssd1 vccd1 vccd1 _13846_/X sky130_fd_sc_hd__o21a_2
XFILLER_90_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_216_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16565_ _18747_/Q _18711_/Q _16565_/S vssd1 vssd1 vccd1 vccd1 _16565_/X sky130_fd_sc_hd__mux2_1
X_13777_ _18657_/Q _13615_/A _13775_/X _13776_/X vssd1 vssd1 vccd1 vccd1 _13777_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_15_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10989_ _14204_/B _09523_/X _10977_/X _10982_/A _18994_/Q vssd1 vssd1 vccd1 vccd1
+ _18998_/D sky130_fd_sc_hd__a32o_1
XFILLER_204_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18304_ _18307_/CLK _18304_/D vssd1 vssd1 vccd1 vccd1 _18304_/Q sky130_fd_sc_hd__dfxtp_1
X_15516_ _15516_/A vssd1 vssd1 vccd1 vccd1 _15516_/X sky130_fd_sc_hd__clkbuf_2
X_12728_ _18094_/Q _18093_/Q _13329_/B vssd1 vssd1 vccd1 vccd1 _12729_/B sky130_fd_sc_hd__or3_1
X_16496_ _16559_/A vssd1 vssd1 vccd1 vccd1 _16496_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_206_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_203_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18235_ _18245_/CLK _18235_/D vssd1 vssd1 vccd1 vccd1 _18235_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15447_ _16962_/A vssd1 vssd1 vccd1 vccd1 _16041_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_175_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12659_ _17931_/Q vssd1 vssd1 vccd1 vccd1 _12662_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_50_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18166_ _18967_/CLK _18166_/D vssd1 vssd1 vccd1 vccd1 _18166_/Q sky130_fd_sc_hd__dfxtp_2
X_15378_ _15982_/A _15393_/B vssd1 vssd1 vccd1 vccd1 _15390_/B sky130_fd_sc_hd__nor2_1
XFILLER_156_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_184_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_156_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17117_ _17197_/A vssd1 vssd1 vccd1 vccd1 _17117_/X sky130_fd_sc_hd__buf_2
XFILLER_50_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14329_ _14275_/X _14326_/X _14328_/X _14270_/X vssd1 vssd1 vccd1 vccd1 _18178_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_89_1366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18097_ _18125_/CLK _18097_/D vssd1 vssd1 vccd1 vccd1 _18097_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_172_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17048_ _17480_/A _17070_/B vssd1 vssd1 vccd1 vccd1 _17056_/B sky130_fd_sc_hd__nor2_1
XFILLER_125_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09870_ _18101_/Q _10627_/B vssd1 vssd1 vccd1 vccd1 _09872_/B sky130_fd_sc_hd__xnor2_1
XFILLER_48_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_225_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18999_ _19000_/CLK _18999_/D vssd1 vssd1 vccd1 vccd1 hold3/A sky130_fd_sc_hd__dfxtp_1
XFILLER_98_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_18 _09209_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_29 _14297_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_227_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_226_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_1304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_199_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_213_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_224_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09304_ _09304_/A _09304_/B _09304_/C _09304_/D vssd1 vssd1 vccd1 vccd1 _09304_/X
+ sky130_fd_sc_hd__and4_1
XFILLER_34_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_221_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09235_ _18917_/Q _18916_/Q _18915_/Q vssd1 vssd1 vccd1 vccd1 _09237_/C sky130_fd_sc_hd__or3_4
XFILLER_139_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_186_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09166_ _18638_/Q _18637_/Q _18636_/Q vssd1 vssd1 vccd1 vccd1 _09170_/A sky130_fd_sc_hd__or3_4
XFILLER_194_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09097_ _18788_/Q _18787_/Q _18786_/Q vssd1 vssd1 vccd1 vccd1 _09098_/D sky130_fd_sc_hd__or3_4
XFILLER_108_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19088__59 vssd1 vssd1 vccd1 vccd1 _19088__59/HI _19196_/A sky130_fd_sc_hd__conb_1
XFILLER_66_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10010_ _10010_/A vssd1 vssd1 vccd1 vccd1 _10010_/X sky130_fd_sc_hd__buf_2
XFILLER_103_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09999_ _09999_/A vssd1 vssd1 vccd1 vccd1 _10086_/A sky130_fd_sc_hd__clkbuf_4
XTAP_5247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_229_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11961_ _12041_/B _11961_/B vssd1 vssd1 vccd1 vccd1 _12026_/B sky130_fd_sc_hd__nor2_2
XTAP_4579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_218_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13700_ _18738_/Q _13642_/X _13582_/A _18744_/Q vssd1 vssd1 vccd1 vccd1 _13700_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_3867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10912_ _10512_/B _10534_/X _10547_/X _10897_/X _10911_/X vssd1 vssd1 vccd1 vccd1
+ _13411_/C sky130_fd_sc_hd__a2111o_1
X_14680_ _18261_/Q _14683_/B _14679_/X _14668_/X vssd1 vssd1 vccd1 vccd1 _18261_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_3878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11892_ _11892_/A _11892_/B _13418_/C vssd1 vssd1 vccd1 vccd1 _11892_/X sky130_fd_sc_hd__or3_1
XFILLER_217_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13631_ _18471_/Q _13531_/A _13630_/X _18447_/Q vssd1 vssd1 vccd1 vccd1 _13631_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_32_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10843_ _13007_/A _10843_/B _10843_/C vssd1 vssd1 vccd1 vccd1 _10843_/X sky130_fd_sc_hd__and3_1
XFILLER_198_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16350_ _16389_/A _16353_/B vssd1 vssd1 vccd1 vccd1 _16350_/Y sky130_fd_sc_hd__nand2_1
X_13562_ _13562_/A vssd1 vssd1 vccd1 vccd1 _13621_/A sky130_fd_sc_hd__buf_6
XFILLER_44_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10774_ _10757_/X _10761_/X _10773_/X vssd1 vssd1 vccd1 vccd1 _10774_/X sky130_fd_sc_hd__a21bo_1
XFILLER_201_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_201_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15301_ _15301_/A _15303_/B vssd1 vssd1 vccd1 vccd1 _15301_/Y sky130_fd_sc_hd__nand2_1
XFILLER_164_1295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12513_ _13153_/A _12513_/B vssd1 vssd1 vccd1 vccd1 _17913_/D sky130_fd_sc_hd__nor2_1
X_16281_ _16285_/B _16277_/X _16280_/Y _16274_/X vssd1 vssd1 vccd1 vccd1 _18640_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_185_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13493_ _13493_/A vssd1 vssd1 vccd1 vccd1 _13493_/X sky130_fd_sc_hd__buf_4
XFILLER_199_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18020_ _18095_/CLK _18020_/D vssd1 vssd1 vccd1 vccd1 _18020_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_60_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15232_ _15232_/A vssd1 vssd1 vccd1 vccd1 _15279_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_12444_ _12446_/A _12444_/B vssd1 vssd1 vccd1 vccd1 _12444_/Y sky130_fd_sc_hd__nand2_1
XFILLER_173_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_138_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15163_ _15169_/B _15161_/X _15162_/X _15143_/X vssd1 vssd1 vccd1 vccd1 _18378_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_197_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12375_ _17894_/Q _12381_/B _12375_/C vssd1 vssd1 vccd1 vccd1 _12375_/Y sky130_fd_sc_hd__nor3_1
XFILLER_5_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14114_ _18938_/Q _13621_/A _13508_/X _18920_/Q vssd1 vssd1 vccd1 vccd1 _14114_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_153_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11326_ _11345_/A _17875_/Q vssd1 vssd1 vccd1 vccd1 _11328_/A sky130_fd_sc_hd__nor2_1
X_15094_ _15118_/A _15094_/B vssd1 vssd1 vccd1 vccd1 _15094_/Y sky130_fd_sc_hd__nand2_1
XFILLER_119_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14045_ _18524_/Q _13642_/X _13841_/A _18530_/Q _14044_/X vssd1 vssd1 vccd1 vccd1
+ _14045_/X sky130_fd_sc_hd__a221o_1
X_18922_ _18959_/CLK _18922_/D vssd1 vssd1 vccd1 vccd1 _18922_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_107_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11257_ _11455_/C _11257_/B _11595_/A vssd1 vssd1 vccd1 vccd1 _11258_/B sky130_fd_sc_hd__or3b_1
XFILLER_79_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_171_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10208_ _10217_/B _10217_/A vssd1 vssd1 vccd1 vccd1 _10210_/B sky130_fd_sc_hd__or2b_1
XFILLER_84_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18853_ _18862_/CLK _18853_/D vssd1 vssd1 vccd1 vccd1 _18853_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_192_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11188_ _11188_/A vssd1 vssd1 vccd1 vccd1 _11210_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_132_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17804_ _17821_/CLK _17804_/D vssd1 vssd1 vccd1 vccd1 _17804_/Q sky130_fd_sc_hd__dfxtp_2
X_10139_ _18119_/Q _10116_/B _09735_/Y vssd1 vssd1 vccd1 vccd1 _10160_/B sky130_fd_sc_hd__a21bo_1
XFILLER_212_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18784_ _18785_/CLK _18784_/D vssd1 vssd1 vccd1 vccd1 _18784_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_94_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15996_ _16193_/A vssd1 vssd1 vccd1 vccd1 _16043_/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_5781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17735_ _17735_/A vssd1 vssd1 vccd1 vccd1 _19011_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_36_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_212_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14947_ _18362_/Q _18326_/Q _14955_/S vssd1 vssd1 vccd1 vccd1 _14947_/X sky130_fd_sc_hd__mux2_1
XFILLER_48_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_224_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_169_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_224_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17666_ _17681_/A _17666_/B vssd1 vssd1 vccd1 vccd1 _17667_/A sky130_fd_sc_hd__and2_1
XFILLER_208_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14878_ _15172_/A _14937_/B vssd1 vssd1 vccd1 vccd1 _14890_/B sky130_fd_sc_hd__nor2_2
XFILLER_62_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINSDIODE2_100 _13848_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_111 _14088_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XINSDIODE2_122 _15233_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_133 _15270_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16617_ _18760_/Q _18724_/Q _16617_/S vssd1 vssd1 vccd1 vccd1 _16617_/X sky130_fd_sc_hd__mux2_1
XFILLER_62_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XINSDIODE2_144 _15589_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13829_ _13829_/A _13829_/B _13829_/C _13829_/D vssd1 vssd1 vccd1 vccd1 _13829_/X
+ sky130_fd_sc_hd__or4_1
XFILLER_50_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17597_ _17610_/A _17597_/B vssd1 vssd1 vccd1 vccd1 _17598_/A sky130_fd_sc_hd__and2_1
XINSDIODE2_155 _18388_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINSDIODE2_166 _18320_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XINSDIODE2_177 _18674_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16548_ _16551_/B _16546_/X _16547_/Y _16539_/X vssd1 vssd1 vccd1 vccd1 _18706_/D
+ sky130_fd_sc_hd__o211a_1
XINSDIODE2_188 _09109_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_199 _10472_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_203_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16479_ _16771_/A _16501_/B vssd1 vssd1 vccd1 vccd1 _16487_/B sky130_fd_sc_hd__nor2_1
XFILLER_176_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09020_ _09022_/A vssd1 vssd1 vccd1 vccd1 _09020_/Y sky130_fd_sc_hd__clkinv_4
X_18218_ _18993_/CLK _18218_/D vssd1 vssd1 vccd1 vccd1 _18218_/Q sky130_fd_sc_hd__dfxtp_1
X_19198_ _19198_/A _08983_/Y vssd1 vssd1 vccd1 vccd1 io_out[36] sky130_fd_sc_hd__ebufn_8
XFILLER_176_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18149_ _18149_/CLK _18149_/D vssd1 vssd1 vccd1 vccd1 _18149_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_145_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09922_ _10294_/A vssd1 vssd1 vccd1 vccd1 _09937_/A sky130_fd_sc_hd__buf_4
XFILLER_160_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_217_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09853_ _09853_/A _09853_/B vssd1 vssd1 vccd1 vccd1 _09853_/Y sky130_fd_sc_hd__nor2_1
XFILLER_24_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_213_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09784_ _09784_/A _09784_/B vssd1 vssd1 vccd1 vccd1 _09787_/A sky130_fd_sc_hd__xnor2_1
XFILLER_230_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_5_31_0_wb_clk_i clkbuf_5_31_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_5_31_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_186_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09218_ _18695_/Q _18694_/Q _18693_/Q vssd1 vssd1 vccd1 vccd1 _09219_/D sky130_fd_sc_hd__or3_4
XFILLER_127_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10490_ _09153_/A _09143_/B _10518_/A vssd1 vssd1 vccd1 vccd1 _10491_/B sky130_fd_sc_hd__mux2_1
XFILLER_10_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09149_ _18713_/Q _18712_/Q _18711_/Q vssd1 vssd1 vccd1 vccd1 _09153_/A sky130_fd_sc_hd__or3_4
XFILLER_107_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12160_ _12157_/Y _12158_/X _12172_/B vssd1 vssd1 vccd1 vccd1 _12160_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_30_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11111_ _11467_/C vssd1 vssd1 vccd1 vccd1 _11654_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_155_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12091_ _12092_/A _12092_/B vssd1 vssd1 vccd1 vccd1 _12091_/X sky130_fd_sc_hd__or2_1
XTAP_5000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11042_ _13344_/A vssd1 vssd1 vccd1 vccd1 _11042_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_110_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_231_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_231_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15850_ _15873_/A _15853_/B vssd1 vssd1 vccd1 vccd1 _15850_/Y sky130_fd_sc_hd__nand2_1
XTAP_5055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14801_ _18326_/Q _18290_/Q _14809_/S vssd1 vssd1 vccd1 vccd1 _14801_/X sky130_fd_sc_hd__mux2_1
XTAP_5099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15781_ _18560_/Q _18524_/Q _15790_/S vssd1 vssd1 vccd1 vccd1 _15781_/X sky130_fd_sc_hd__mux2_1
XTAP_4365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12993_ _12990_/A _13007_/B _12992_/X _12972_/X vssd1 vssd1 vccd1 vccd1 _17978_/D
+ sky130_fd_sc_hd__a211o_1
XFILLER_92_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17520_ _18979_/Q _18943_/Q _17533_/S vssd1 vssd1 vccd1 vccd1 _17520_/X sky130_fd_sc_hd__mux2_1
XFILLER_91_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14732_ _15172_/A _14790_/B vssd1 vssd1 vccd1 vccd1 _14742_/B sky130_fd_sc_hd__nor2_2
XFILLER_29_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_217_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11944_ _11944_/A _12025_/B _13426_/A _11999_/C vssd1 vssd1 vccd1 vccd1 _11944_/X
+ sky130_fd_sc_hd__or4_2
XFILLER_91_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17451_ _17519_/A vssd1 vssd1 vccd1 vccd1 _17467_/S sky130_fd_sc_hd__clkbuf_2
XTAP_2963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14663_ _16932_/A vssd1 vssd1 vccd1 vccd1 _16935_/A sky130_fd_sc_hd__buf_4
XFILLER_33_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11875_ _11868_/B _11860_/B _11869_/Y vssd1 vssd1 vccd1 vccd1 _11875_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_44_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16402_ _16447_/A _16407_/B vssd1 vssd1 vccd1 vccd1 _16402_/Y sky130_fd_sc_hd__nand2_1
XFILLER_44_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_220_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13614_ _13738_/A vssd1 vssd1 vccd1 vccd1 _13615_/A sky130_fd_sc_hd__buf_2
X_10826_ _10826_/A _10877_/B vssd1 vssd1 vccd1 vccd1 _10826_/X sky130_fd_sc_hd__or2_1
X_17382_ _18944_/Q _18908_/Q _17386_/S vssd1 vssd1 vccd1 vccd1 _17382_/X sky130_fd_sc_hd__mux2_1
XFILLER_207_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14594_ _16862_/A vssd1 vssd1 vccd1 vccd1 _15197_/A sky130_fd_sc_hd__buf_8
XFILLER_38_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16333_ _16371_/A _16773_/B _16333_/C vssd1 vssd1 vccd1 vccd1 _16333_/X sky130_fd_sc_hd__or3_1
X_13545_ _14016_/A vssd1 vssd1 vccd1 vccd1 _13546_/A sky130_fd_sc_hd__buf_8
X_10757_ _10757_/A _10757_/B _10757_/C vssd1 vssd1 vccd1 vccd1 _10757_/X sky130_fd_sc_hd__or3_1
XFILLER_9_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16264_ _18673_/Q _18637_/Q _16271_/S vssd1 vssd1 vccd1 vccd1 _16264_/X sky130_fd_sc_hd__mux2_1
X_13476_ _17845_/Q _13459_/X _12184_/X vssd1 vssd1 vccd1 vccd1 _18161_/D sky130_fd_sc_hd__o21a_1
XFILLER_12_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10688_ _09277_/A _09277_/B _09277_/C _09277_/D _10695_/A _10764_/A vssd1 vssd1 vccd1
+ vccd1 _10689_/C sky130_fd_sc_hd__mux4_2
XFILLER_127_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_1330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18003_ _18997_/CLK _18003_/D vssd1 vssd1 vccd1 vccd1 _18003_/Q sky130_fd_sc_hd__dfxtp_1
X_15215_ _18391_/Q _15216_/B _15214_/Y _15208_/X vssd1 vssd1 vccd1 vccd1 _18391_/D
+ sky130_fd_sc_hd__o211a_1
X_12427_ _12427_/A vssd1 vssd1 vccd1 vccd1 _12429_/A sky130_fd_sc_hd__inv_2
X_16195_ _16248_/A _16785_/B _16208_/C vssd1 vssd1 vccd1 vccd1 _16195_/X sky130_fd_sc_hd__or3_1
XFILLER_154_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15146_ _15211_/A vssd1 vssd1 vccd1 vccd1 _15279_/C sky130_fd_sc_hd__clkbuf_2
X_12358_ _12486_/B _12358_/B vssd1 vssd1 vccd1 vccd1 _12495_/A sky130_fd_sc_hd__nand2_1
XFILLER_114_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11309_ _11735_/B _11617_/A _11305_/X _11308_/Y vssd1 vssd1 vccd1 vccd1 _11310_/C
+ sky130_fd_sc_hd__o31a_1
XFILLER_99_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15077_ _15082_/B _15075_/X _15076_/X _15066_/X vssd1 vssd1 vccd1 vccd1 _18357_/D
+ sky130_fd_sc_hd__o211a_1
X_12289_ _12289_/A _12304_/B vssd1 vssd1 vccd1 vccd1 _12300_/A sky130_fd_sc_hd__nor2_1
X_14028_ _18248_/Q _13877_/X _13515_/A _18242_/Q vssd1 vssd1 vccd1 vccd1 _14028_/X
+ sky130_fd_sc_hd__a22o_1
X_18905_ _18908_/CLK _18905_/D vssd1 vssd1 vccd1 vccd1 _18905_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_45_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_136_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18836_ _18871_/CLK _18836_/D vssd1 vssd1 vccd1 vccd1 _18836_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_45_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_212_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18767_ _18773_/CLK _18767_/D vssd1 vssd1 vccd1 vccd1 _18767_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15979_ _18571_/Q _15980_/B _15978_/Y _15972_/X vssd1 vssd1 vccd1 vccd1 _18571_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_110_1323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_208_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17718_ _17718_/A vssd1 vssd1 vccd1 vccd1 _19003_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_224_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18698_ _18732_/CLK _18698_/D vssd1 vssd1 vccd1 vccd1 _18698_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_63_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_1367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17649_ _17674_/A _17663_/B vssd1 vssd1 vccd1 vccd1 _17649_/Y sky130_fd_sc_hd__nor2_1
XFILLER_91_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_177_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_211_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_189_wb_clk_i clkbuf_5_9_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18163_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_56_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_182_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_1274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_118_wb_clk_i clkbuf_5_28_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18506_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_143_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_192_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09003_ _09003_/A vssd1 vssd1 vccd1 vccd1 _09003_/Y sky130_fd_sc_hd__inv_2
XFILLER_178_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_219_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_219_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19058__29 vssd1 vssd1 vccd1 vccd1 _19058__29/HI _19152_/A sky130_fd_sc_hd__conb_1
XFILLER_63_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09905_ _09905_/A vssd1 vssd1 vccd1 vccd1 _09905_/X sky130_fd_sc_hd__buf_4
XFILLER_154_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_219_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09836_ _18100_/Q vssd1 vssd1 vccd1 vccd1 _13348_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_150_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_189_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09767_ _18123_/Q vssd1 vssd1 vccd1 vccd1 _09774_/A sky130_fd_sc_hd__inv_2
XFILLER_100_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09698_ _18266_/Q _18265_/Q _18264_/Q vssd1 vssd1 vccd1 vccd1 _09698_/X sky130_fd_sc_hd__or3_4
XFILLER_73_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_215_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_214_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_187_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11660_ _11653_/Y _11665_/B _11705_/D vssd1 vssd1 vccd1 vccd1 _11683_/B sky130_fd_sc_hd__a21o_1
XPHY_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_230_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10611_ _18129_/Q _10611_/B vssd1 vssd1 vccd1 vccd1 _10612_/B sky130_fd_sc_hd__nor2_1
XFILLER_186_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11591_ _11268_/Y _11591_/B vssd1 vssd1 vccd1 vccd1 _11592_/D sky130_fd_sc_hd__and2b_1
XFILLER_122_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_195_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13330_ _18094_/Q _13329_/X _11891_/X vssd1 vssd1 vccd1 vccd1 _13330_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_22_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_195_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10542_ _10542_/A vssd1 vssd1 vccd1 vccd1 _10542_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_109_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13261_ _13261_/A vssd1 vssd1 vccd1 vccd1 _18083_/D sky130_fd_sc_hd__clkbuf_1
X_10473_ _09248_/A _09243_/A _09253_/B _10097_/A _10462_/X _10450_/S vssd1 vssd1 vccd1
+ vccd1 _10474_/B sky130_fd_sc_hd__mux4_1
XFILLER_202_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15000_ _15064_/A vssd1 vssd1 vccd1 vccd1 _15134_/B sky130_fd_sc_hd__buf_2
X_12212_ _11691_/Y _12210_/A _12209_/X _12239_/C _12147_/X vssd1 vssd1 vccd1 vccd1
+ _17852_/D sky130_fd_sc_hd__o2111a_1
XFILLER_6_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13192_ _13192_/A vssd1 vssd1 vccd1 vccd1 _18052_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_123_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12143_ _13458_/A vssd1 vssd1 vccd1 vccd1 _12183_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_150_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16951_ _16957_/B _16947_/X _16950_/X _16940_/X vssd1 vssd1 vccd1 vccd1 _18801_/D
+ sky130_fd_sc_hd__o211a_1
X_12074_ _12074_/A vssd1 vssd1 vccd1 vccd1 _12975_/A sky130_fd_sc_hd__buf_4
XFILLER_111_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15902_ _15900_/B _15899_/X _15900_/Y _15901_/X vssd1 vssd1 vccd1 vccd1 _18554_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_49_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11025_ _11044_/A _11025_/B vssd1 vssd1 vccd1 vccd1 _11026_/A sky130_fd_sc_hd__nand2_1
XFILLER_110_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16882_ _16882_/A _16884_/B vssd1 vssd1 vccd1 vccd1 _16882_/Y sky130_fd_sc_hd__nand2_1
XFILLER_133_1367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18621_ _18623_/CLK _18621_/D vssd1 vssd1 vccd1 vccd1 _18621_/Q sky130_fd_sc_hd__dfxtp_2
X_15833_ _15857_/A _15984_/B _15870_/C vssd1 vssd1 vccd1 vccd1 _15833_/X sky130_fd_sc_hd__or3_1
XTAP_4140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19072__43 vssd1 vssd1 vccd1 vccd1 _19072__43/HI _19166_/A sky130_fd_sc_hd__conb_1
XFILLER_49_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18552_ _18553_/CLK _18552_/D vssd1 vssd1 vccd1 vccd1 _18552_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_4184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15764_ _18519_/Q _15769_/B _15762_/X _15763_/X vssd1 vssd1 vccd1 vccd1 _18519_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_4195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12976_ _12976_/A _12976_/B vssd1 vssd1 vccd1 vccd1 _12976_/X sky130_fd_sc_hd__or2_1
XFILLER_92_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_206_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17503_ _17503_/A _17536_/B vssd1 vssd1 vccd1 vccd1 _17512_/B sky130_fd_sc_hd__nor2_2
XTAP_3483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14715_ _14753_/A _14715_/B vssd1 vssd1 vccd1 vccd1 _14715_/Y sky130_fd_sc_hd__nand2_1
XFILLER_18_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18483_ _18506_/CLK _18483_/D vssd1 vssd1 vccd1 vccd1 _18483_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11927_ _11927_/A vssd1 vssd1 vccd1 vccd1 _11932_/A sky130_fd_sc_hd__clkbuf_2
X_15695_ _15694_/B _15693_/X _15694_/Y _15681_/X vssd1 vssd1 vccd1 vccd1 _18503_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_2760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17434_ _17472_/A vssd1 vssd1 vccd1 vccd1 _17491_/B sky130_fd_sc_hd__buf_2
XFILLER_162_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14646_ _14683_/A _14646_/B vssd1 vssd1 vccd1 vccd1 _14646_/Y sky130_fd_sc_hd__nand2_1
XFILLER_33_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11858_ _11778_/X _11856_/X _11857_/Y _11809_/X vssd1 vssd1 vccd1 vccd1 _11858_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_33_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17365_ _17376_/A _17506_/B _17376_/C vssd1 vssd1 vccd1 vccd1 _17365_/X sky130_fd_sc_hd__or3_1
X_10809_ _10809_/A _10809_/B vssd1 vssd1 vccd1 vccd1 _10809_/X sky130_fd_sc_hd__or2_1
XFILLER_203_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11789_ _11789_/A _13429_/A vssd1 vssd1 vccd1 vccd1 _11789_/Y sky130_fd_sc_hd__nand2_1
X_14577_ _18171_/Q _18172_/Q vssd1 vssd1 vccd1 vccd1 _14685_/B sky130_fd_sc_hd__or2b_1
XFILLER_159_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_211_wb_clk_i clkbuf_5_12_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17821_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_16316_ _18686_/Q _18650_/Q _16324_/S vssd1 vssd1 vccd1 vccd1 _16316_/X sky130_fd_sc_hd__mux2_1
XFILLER_192_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13528_ _13670_/A vssd1 vssd1 vccd1 vccd1 _13529_/A sky130_fd_sc_hd__buf_4
XFILLER_119_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_1338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17296_ _17318_/A _17437_/B _17318_/C vssd1 vssd1 vccd1 vccd1 _17296_/X sky130_fd_sc_hd__or3_1
XFILLER_201_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19035_ _19035_/CLK _19035_/D vssd1 vssd1 vccd1 vccd1 _19035_/Q sky130_fd_sc_hd__dfxtp_1
X_16247_ _18669_/Q _18633_/Q _16250_/S vssd1 vssd1 vccd1 vccd1 _16247_/X sky130_fd_sc_hd__mux2_1
XFILLER_173_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13459_ _13465_/A vssd1 vssd1 vccd1 vccd1 _13459_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_63_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16178_ _16771_/A _16205_/B vssd1 vssd1 vccd1 vccd1 _16188_/B sky130_fd_sc_hd__nor2_2
XFILLER_142_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15129_ _15132_/B _15126_/X _15128_/Y _15123_/X vssd1 vssd1 vccd1 vccd1 _18370_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_142_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_229_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09621_ _18104_/Q vssd1 vssd1 vccd1 vccd1 _10204_/A sky130_fd_sc_hd__buf_2
X_18819_ _18826_/CLK _18819_/D vssd1 vssd1 vccd1 vccd1 _18819_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_56_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09552_ _09565_/A vssd1 vssd1 vccd1 vccd1 _10123_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_23_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09483_ _09483_/A vssd1 vssd1 vccd1 vccd1 _18148_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_64_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_212_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_177_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_211_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_139_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_191_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_86_wb_clk_i _18144_/CLK vssd1 vssd1 vccd1 vccd1 _18590_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_219_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_191_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_15_wb_clk_i clkbuf_5_4_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18893_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_8_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_219_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09819_ _10403_/A vssd1 vssd1 vccd1 vccd1 _12133_/A sky130_fd_sc_hd__buf_2
XFILLER_115_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_219_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12830_ _12699_/Y _12913_/A _12542_/B _12846_/A vssd1 vssd1 vccd1 vccd1 _12830_/X
+ sky130_fd_sc_hd__a2bb2o_1
XTAP_2012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12761_ _13318_/C _12747_/Y _12760_/X vssd1 vssd1 vccd1 vccd1 _12761_/X sky130_fd_sc_hd__o21a_1
XTAP_2056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14500_ _18224_/Q _14502_/B vssd1 vssd1 vccd1 vccd1 _14501_/A sky130_fd_sc_hd__and2_1
XTAP_1333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11712_ _13452_/A _11286_/X _11681_/C vssd1 vssd1 vccd1 vccd1 _11712_/X sky130_fd_sc_hd__o21a_1
XTAP_1344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15480_ _18486_/Q _18450_/Q _15494_/S vssd1 vssd1 vccd1 vccd1 _15480_/X sky130_fd_sc_hd__mux2_1
XFILLER_15_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12692_ _12707_/A _12662_/A _12688_/Y vssd1 vssd1 vccd1 vccd1 _12693_/B sky130_fd_sc_hd__o21ai_1
XFILLER_230_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11643_ _17860_/Q vssd1 vssd1 vccd1 vccd1 _11671_/B sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_1388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14431_ _14422_/X _09500_/B _14423_/X vssd1 vssd1 vccd1 vccd1 _14431_/X sky130_fd_sc_hd__a21o_1
XTAP_1399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17150_ _17156_/B _17147_/X _17149_/X _17140_/X vssd1 vssd1 vccd1 vccd1 _18849_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_35_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11574_ _11253_/A _11495_/B _11547_/Y _11366_/A _11573_/Y vssd1 vssd1 vccd1 vccd1
+ _11574_/X sky130_fd_sc_hd__o2111a_1
X_14362_ _17944_/Q _14272_/X _14361_/X _12972_/X vssd1 vssd1 vccd1 vccd1 _18184_/D
+ sky130_fd_sc_hd__a211o_1
XFILLER_7_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_168_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16101_ _18636_/Q _18600_/Q _16113_/S vssd1 vssd1 vccd1 vccd1 _16101_/X sky130_fd_sc_hd__mux2_1
XFILLER_168_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10525_ _10523_/X _10524_/X _10935_/S vssd1 vssd1 vccd1 vccd1 _10525_/X sky130_fd_sc_hd__mux2_2
XFILLER_155_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13313_ _13314_/A vssd1 vssd1 vccd1 vccd1 _13313_/X sky130_fd_sc_hd__clkbuf_2
X_17081_ _17080_/B _17079_/X _17080_/Y _17076_/X vssd1 vssd1 vccd1 vccd1 _18833_/D
+ sky130_fd_sc_hd__o211a_1
X_14293_ _14293_/A _14293_/B vssd1 vssd1 vccd1 vccd1 _14294_/B sky130_fd_sc_hd__nor2_1
XFILLER_6_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_1300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_196_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16032_ _16043_/A _16032_/B _16043_/C vssd1 vssd1 vccd1 vccd1 _16032_/X sky130_fd_sc_hd__or3_1
XFILLER_7_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13244_ _13244_/A _18077_/Q vssd1 vssd1 vccd1 vccd1 _13245_/A sky130_fd_sc_hd__and2_1
XFILLER_143_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10456_ _10456_/A _12031_/A vssd1 vssd1 vccd1 vccd1 _10512_/B sky130_fd_sc_hd__nor2_2
XFILLER_108_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_182_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13175_ _13175_/A _18046_/Q vssd1 vssd1 vccd1 vccd1 _13176_/A sky130_fd_sc_hd__and2_1
XFILLER_83_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10387_ _09344_/C _09344_/D _09354_/D _09349_/D _09972_/B _09959_/A vssd1 vssd1 vccd1
+ vccd1 _10388_/B sky130_fd_sc_hd__mux4_2
XFILLER_124_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12126_ _12126_/A _12126_/B vssd1 vssd1 vccd1 vccd1 _12127_/D sky130_fd_sc_hd__xor2_1
XFILLER_124_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17983_ _18044_/CLK _17983_/D vssd1 vssd1 vccd1 vccd1 _17983_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_81_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16934_ _18834_/Q _18798_/Q _16947_/S vssd1 vssd1 vccd1 vccd1 _16934_/X sky130_fd_sc_hd__mux2_1
XFILLER_46_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12057_ _13518_/B vssd1 vssd1 vccd1 vccd1 _13526_/B sky130_fd_sc_hd__inv_2
XFILLER_78_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11008_ _17813_/Q _11201_/A _17811_/Q _11196_/B vssd1 vssd1 vccd1 vccd1 _11011_/C
+ sky130_fd_sc_hd__nand4_1
XFILLER_77_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16865_ _16865_/A vssd1 vssd1 vccd1 vccd1 _17460_/B sky130_fd_sc_hd__buf_6
XFILLER_37_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_226_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_225_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18604_ _18607_/CLK _18604_/D vssd1 vssd1 vccd1 vccd1 _18604_/Q sky130_fd_sc_hd__dfxtp_2
X_15816_ _15818_/B _15814_/X _15815_/Y _15803_/X vssd1 vssd1 vccd1 vccd1 _18532_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_168_1238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16796_ _16796_/A _16796_/B _16796_/C vssd1 vssd1 vccd1 vccd1 _16796_/X sky130_fd_sc_hd__or3_1
XFILLER_225_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18535_ _18546_/CLK _18535_/D vssd1 vssd1 vccd1 vccd1 _18535_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_209_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15747_ _15869_/A vssd1 vssd1 vccd1 vccd1 _15799_/A sky130_fd_sc_hd__clkbuf_2
XTAP_3280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12959_ _12969_/A _12959_/B vssd1 vssd1 vccd1 vccd1 _12961_/B sky130_fd_sc_hd__nor2_1
XFILLER_46_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_221_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18466_ _18467_/CLK _18466_/D vssd1 vssd1 vccd1 vccd1 _18466_/Q sky130_fd_sc_hd__dfxtp_2
X_15678_ _15678_/A _16128_/B _15724_/C vssd1 vssd1 vccd1 vccd1 _15678_/X sky130_fd_sc_hd__or3_1
XTAP_2590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17417_ _17453_/A _17419_/B vssd1 vssd1 vccd1 vccd1 _17417_/Y sky130_fd_sc_hd__nand2_1
X_14629_ _14668_/A vssd1 vssd1 vccd1 vccd1 _14629_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_53_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_221_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18397_ _18398_/CLK _18397_/D vssd1 vssd1 vccd1 vccd1 _18397_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_33_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_221_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17348_ _17468_/A vssd1 vssd1 vccd1 vccd1 _17395_/A sky130_fd_sc_hd__buf_2
XFILLER_179_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17279_ _17390_/A vssd1 vssd1 vccd1 vccd1 _17370_/A sky130_fd_sc_hd__buf_2
XFILLER_179_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_179_1367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19018_ _19019_/CLK _19018_/D vssd1 vssd1 vccd1 vccd1 _19018_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_134_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_146_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_3_0_0_wb_clk_i clkbuf_3_1_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_4_1_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_138_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_216_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08983_ _08985_/A vssd1 vssd1 vccd1 vccd1 _08983_/Y sky130_fd_sc_hd__inv_2
XFILLER_25_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_229_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_217_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_1305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09604_ _13005_/A vssd1 vssd1 vccd1 vccd1 _10155_/C sky130_fd_sc_hd__inv_2
XFILLER_112_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09535_ _18103_/Q _09535_/B vssd1 vssd1 vccd1 vccd1 _10114_/B sky130_fd_sc_hd__xnor2_4
XFILLER_227_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_133_wb_clk_i clkbuf_5_24_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18408_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_225_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09466_ _09475_/A _09466_/B vssd1 vssd1 vccd1 vccd1 _09467_/B sky130_fd_sc_hd__and2_1
XFILLER_24_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_227_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_212_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_196_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09397_ _09397_/A _09397_/B _09397_/C _09397_/D vssd1 vssd1 vccd1 vccd1 _09403_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_36_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10310_ _10291_/X _10307_/X _10309_/X _10370_/S vssd1 vssd1 vccd1 vccd1 _10310_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_192_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_180_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11290_ _11354_/B _11289_/X _11681_/D vssd1 vssd1 vccd1 vccd1 _11303_/A sky130_fd_sc_hd__mux2_1
XFILLER_3_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10241_ _10521_/A vssd1 vssd1 vccd1 vccd1 _10561_/S sky130_fd_sc_hd__buf_2
XFILLER_152_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_133_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10172_ _10172_/A _10172_/B _10172_/C vssd1 vssd1 vccd1 vccd1 _12053_/B sky130_fd_sc_hd__nand3_1
XFILLER_191_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14980_ _14980_/A vssd1 vssd1 vccd1 vccd1 _14980_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_43_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13931_ _18265_/Q _13714_/X _13698_/A _18256_/Q _13930_/X vssd1 vssd1 vccd1 vccd1
+ _13931_/X sky130_fd_sc_hd__a221o_1
XFILLER_130_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16650_ _16794_/A _16650_/B vssd1 vssd1 vccd1 vccd1 _16658_/B sky130_fd_sc_hd__nor2_2
XFILLER_170_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19042__13 vssd1 vssd1 vccd1 vccd1 _19042__13/HI _19136_/A sky130_fd_sc_hd__conb_1
X_13862_ _18811_/Q _13508_/A _13861_/X _18835_/Q vssd1 vssd1 vccd1 vccd1 _13862_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_47_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15601_ _18517_/Q _18481_/Q _15604_/S vssd1 vssd1 vccd1 vccd1 _15601_/X sky130_fd_sc_hd__mux2_1
XFILLER_170_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12813_ _12813_/A _12813_/B _12813_/C _12813_/D vssd1 vssd1 vccd1 vccd1 _12813_/X
+ sky130_fd_sc_hd__or4_1
XFILLER_216_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16581_ _16659_/A vssd1 vssd1 vccd1 vccd1 _16581_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_28_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13793_ _18270_/Q _13735_/X _13764_/X _18294_/Q vssd1 vssd1 vccd1 vccd1 _13793_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_128_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18320_ _18324_/CLK _18320_/D vssd1 vssd1 vccd1 vccd1 _18320_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_43_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15532_ _15566_/A _15534_/B vssd1 vssd1 vccd1 vccd1 _15532_/Y sky130_fd_sc_hd__nand2_1
XFILLER_188_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12744_ _18089_/Q _13318_/A vssd1 vssd1 vccd1 vccd1 _12748_/B sky130_fd_sc_hd__or2_1
XFILLER_215_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_231_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18251_ _18251_/CLK _18251_/D vssd1 vssd1 vccd1 vccd1 _18251_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15463_ _15607_/B _15463_/B _15607_/C vssd1 vssd1 vccd1 vccd1 _17265_/A sky130_fd_sc_hd__nand3b_4
XFILLER_230_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12675_ _17933_/Q vssd1 vssd1 vccd1 vccd1 _12676_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_231_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_204_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17202_ _17491_/A _17202_/B vssd1 vssd1 vccd1 vccd1 _17213_/B sky130_fd_sc_hd__nor2_1
X_14414_ _14414_/A _14414_/B vssd1 vssd1 vccd1 vccd1 _14414_/Y sky130_fd_sc_hd__nor2_1
XFILLER_187_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11626_ _11602_/B _11623_/Y _12235_/A _11625_/X _11689_/A vssd1 vssd1 vccd1 vccd1
+ _11626_/X sky130_fd_sc_hd__a32o_1
X_18182_ _18182_/CLK _18182_/D vssd1 vssd1 vccd1 vccd1 _18182_/Q sky130_fd_sc_hd__dfxtp_4
X_15394_ _15415_/A vssd1 vssd1 vccd1 vccd1 _15412_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_156_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17133_ _17247_/A vssd1 vssd1 vccd1 vccd1 _17226_/A sky130_fd_sc_hd__clkbuf_2
X_14345_ _18180_/Q vssd1 vssd1 vccd1 vccd1 _17119_/A sky130_fd_sc_hd__clkbuf_2
X_11557_ _17866_/Q _17865_/Q vssd1 vssd1 vccd1 vccd1 _12269_/A sky130_fd_sc_hd__and2_1
XFILLER_7_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10508_ _09114_/C _10350_/A _10509_/S vssd1 vssd1 vccd1 vccd1 _10508_/X sky130_fd_sc_hd__mux2_1
X_17064_ _18865_/Q _18829_/Q _17074_/S vssd1 vssd1 vccd1 vccd1 _17064_/X sky130_fd_sc_hd__mux2_1
XFILLER_183_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11488_ _11488_/A _11488_/B vssd1 vssd1 vccd1 vccd1 _11488_/Y sky130_fd_sc_hd__nor2_1
X_14276_ _14187_/A _12066_/A _12099_/A _14237_/A _19000_/Q vssd1 vssd1 vccd1 vccd1
+ _14276_/X sky130_fd_sc_hd__a221o_1
XFILLER_155_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16015_ _18617_/Q _18581_/Q _16031_/S vssd1 vssd1 vccd1 vccd1 _16015_/X sky130_fd_sc_hd__mux2_1
X_13227_ _13233_/A _18069_/Q vssd1 vssd1 vccd1 vccd1 _13228_/A sky130_fd_sc_hd__and2_1
X_10439_ _10424_/X _10436_/Y _10547_/B vssd1 vssd1 vccd1 vccd1 _10439_/X sky130_fd_sc_hd__a21bo_1
XFILLER_83_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13158_ _13164_/A _18038_/Q vssd1 vssd1 vccd1 vccd1 _13159_/A sky130_fd_sc_hd__and2_1
XFILLER_98_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12109_ _09842_/B _12109_/B vssd1 vssd1 vccd1 vccd1 _12109_/X sky130_fd_sc_hd__and2b_1
XFILLER_111_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13089_ _13089_/A vssd1 vssd1 vccd1 vccd1 _18006_/D sky130_fd_sc_hd__clkbuf_1
X_17966_ _17969_/CLK _17966_/D vssd1 vssd1 vccd1 vccd1 _17966_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_100_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16917_ _16999_/A vssd1 vssd1 vccd1 vccd1 _16917_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_120_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17897_ _17919_/CLK _17897_/D vssd1 vssd1 vccd1 vccd1 _17897_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_226_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_225_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16848_ _16871_/A vssd1 vssd1 vccd1 vccd1 _16848_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_226_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_168_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16779_ _16815_/A _16779_/B vssd1 vssd1 vccd1 vccd1 _16779_/Y sky130_fd_sc_hd__nand2_1
XFILLER_213_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09320_ _09320_/A _09320_/B _09320_/C vssd1 vssd1 vccd1 vccd1 _09321_/A sky130_fd_sc_hd__nand3_1
X_18518_ _18553_/CLK _18518_/D vssd1 vssd1 vccd1 vccd1 _18518_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_178_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_1298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09251_ _18902_/Q _18901_/Q _18900_/Q vssd1 vssd1 vccd1 vccd1 _09253_/C sky130_fd_sc_hd__or3_4
X_18449_ _18473_/CLK _18449_/D vssd1 vssd1 vccd1 vccd1 _18449_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_22_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_221_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09182_ _18599_/Q _18598_/Q _18597_/Q vssd1 vssd1 vccd1 vccd1 _09186_/A sky130_fd_sc_hd__or3_2
XFILLER_119_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_175_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08966_ _08966_/A vssd1 vssd1 vccd1 vccd1 _08966_/Y sky130_fd_sc_hd__inv_2
XFILLER_103_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_229_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_217_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_217_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_227_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09518_ _09517_/Y _09518_/B vssd1 vssd1 vccd1 vccd1 _09518_/X sky130_fd_sc_hd__and2b_1
XFILLER_25_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10790_ _10805_/A _10790_/B _10790_/C vssd1 vssd1 vccd1 vccd1 _10790_/X sky130_fd_sc_hd__and3_1
XPHY_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_223_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_197_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_169_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09449_ _09255_/A _09254_/Y _09440_/Y _09448_/Y vssd1 vssd1 vccd1 vccd1 _09463_/A
+ sky130_fd_sc_hd__o211ai_2
XPHY_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_212_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_212_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12460_ _12460_/A vssd1 vssd1 vccd1 vccd1 _17904_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_12_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_228_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_200_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11411_ _11466_/B _11467_/C _11307_/B _11467_/D vssd1 vssd1 vccd1 vccd1 _11594_/A
+ sky130_fd_sc_hd__o31a_1
XFILLER_165_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12391_ _12401_/B vssd1 vssd1 vccd1 vccd1 _12394_/B sky130_fd_sc_hd__inv_2
XFILLER_166_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14130_ _18284_/Q _13877_/X _13842_/A _18278_/Q _14129_/X vssd1 vssd1 vccd1 vccd1
+ _14130_/X sky130_fd_sc_hd__a221o_1
XFILLER_125_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11342_ _11329_/Y _11332_/X _11339_/Y _11645_/A vssd1 vssd1 vccd1 vccd1 _11342_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_193_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_197_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_30_wb_clk_i clkbuf_5_7_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18931_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_4_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14061_ _18395_/Q _13523_/A _13537_/A _18377_/Q vssd1 vssd1 vccd1 vccd1 _14061_/X
+ sky130_fd_sc_hd__a22o_1
X_11273_ _11926_/B _11297_/B vssd1 vssd1 vccd1 vccd1 _11832_/B sky130_fd_sc_hd__or2_1
XFILLER_10_1366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13012_ _13009_/A _12991_/X _13010_/X _13011_/X vssd1 vssd1 vccd1 vccd1 _17982_/D
+ sky130_fd_sc_hd__o211a_1
X_10224_ _10475_/A vssd1 vssd1 vccd1 vccd1 _10555_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_152_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17820_ _17821_/CLK _17820_/D vssd1 vssd1 vccd1 vccd1 _17820_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_79_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10155_ _10155_/A _13389_/A _10155_/C vssd1 vssd1 vccd1 vccd1 _10155_/X sky130_fd_sc_hd__and3_1
XTAP_5930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17751_ _17751_/A vssd1 vssd1 vccd1 vccd1 _19018_/D sky130_fd_sc_hd__clkbuf_1
XTAP_5963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14963_ _15255_/A _14985_/B vssd1 vssd1 vccd1 vccd1 _14971_/B sky130_fd_sc_hd__nor2_1
X_10086_ _10086_/A _10086_/B vssd1 vssd1 vccd1 vccd1 _10086_/Y sky130_fd_sc_hd__nand2_1
XTAP_5974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16702_ _18780_/Q _18744_/Q _16715_/S vssd1 vssd1 vccd1 vccd1 _16702_/X sky130_fd_sc_hd__mux2_1
XFILLER_75_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13914_ _13693_/Y _13897_/X _13905_/X _13913_/X vssd1 vssd1 vccd1 vccd1 _13914_/X
+ sky130_fd_sc_hd__a211o_2
X_17682_ _17682_/A vssd1 vssd1 vccd1 vccd1 _18982_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_78_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14894_ _14919_/A _15186_/B _14906_/C vssd1 vssd1 vccd1 vccd1 _14894_/X sky130_fd_sc_hd__or3_1
XFILLER_35_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_223_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16633_ _18764_/Q _18728_/Q _16637_/S vssd1 vssd1 vccd1 vccd1 _16633_/X sky130_fd_sc_hd__mux2_1
XFILLER_63_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_223_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13845_ _18667_/Q _13508_/X _13839_/X _13844_/X vssd1 vssd1 vccd1 vccd1 _13845_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_74_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_188_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16564_ _16714_/A _16602_/B vssd1 vssd1 vccd1 vccd1 _16575_/B sky130_fd_sc_hd__nor2_1
X_13776_ _18645_/Q _13723_/X _13743_/X _18627_/Q vssd1 vssd1 vccd1 vccd1 _13776_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_50_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10988_ _18998_/Q vssd1 vssd1 vccd1 vccd1 _14204_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_206_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18303_ _18307_/CLK _18303_/D vssd1 vssd1 vccd1 vccd1 _18303_/Q sky130_fd_sc_hd__dfxtp_1
X_15515_ _15551_/A _15964_/B _15515_/C vssd1 vssd1 vccd1 vccd1 _15515_/X sky130_fd_sc_hd__or3_1
X_12727_ _18092_/Q _13322_/B vssd1 vssd1 vccd1 vccd1 _13329_/B sky130_fd_sc_hd__or2_1
X_16495_ _16507_/A _16499_/B vssd1 vssd1 vccd1 vccd1 _16495_/Y sky130_fd_sc_hd__nand2_1
XFILLER_230_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18234_ _18263_/CLK _18234_/D vssd1 vssd1 vccd1 vccd1 _18234_/Q sky130_fd_sc_hd__dfxtp_1
X_15446_ _15445_/B _15444_/X _15445_/Y _15428_/X vssd1 vssd1 vccd1 vccd1 _18443_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_31_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12658_ _17930_/Q _12635_/X _12656_/Y _12657_/X _12621_/X vssd1 vssd1 vccd1 vccd1
+ _17930_/D sky130_fd_sc_hd__a221o_1
XFILLER_141_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11609_ _11609_/A _11617_/B _11786_/B vssd1 vssd1 vccd1 vccd1 _11609_/X sky130_fd_sc_hd__or3_2
X_18165_ _19021_/CLK _18165_/D vssd1 vssd1 vccd1 vccd1 hold2/A sky130_fd_sc_hd__dfxtp_1
X_15377_ _16889_/A vssd1 vssd1 vccd1 vccd1 _15982_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_129_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12589_ _12589_/A _12589_/B vssd1 vssd1 vccd1 vccd1 _12590_/B sky130_fd_sc_hd__nand2_1
XFILLER_157_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17116_ _17323_/A vssd1 vssd1 vccd1 vccd1 _17197_/A sky130_fd_sc_hd__buf_2
XFILLER_7_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14328_ _14299_/X _14282_/X _14283_/X _14300_/X _16512_/C vssd1 vssd1 vccd1 vccd1
+ _14328_/X sky130_fd_sc_hd__a311o_1
XFILLER_209_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18096_ _19028_/CLK _18096_/D vssd1 vssd1 vccd1 vccd1 _18096_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_183_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17047_ _18824_/Q _17046_/B _17046_/Y _17040_/X vssd1 vssd1 vccd1 vccd1 _18824_/D
+ sky130_fd_sc_hd__o211a_1
X_14259_ _12039_/A _14205_/X _14258_/X vssd1 vssd1 vccd1 vccd1 _14259_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_217_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18998_ _19000_/CLK _18998_/D vssd1 vssd1 vccd1 vccd1 _18998_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_19 _09214_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_1215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17949_ _17954_/CLK _17949_/D vssd1 vssd1 vccd1 vccd1 _17949_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_85_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_226_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_226_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_213_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_198_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_5_21_0_wb_clk_i clkbuf_5_21_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_5_21_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_213_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_181_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09303_ _18512_/Q _18511_/Q _18510_/Q vssd1 vssd1 vccd1 vccd1 _09304_/D sky130_fd_sc_hd__or3_4
XFILLER_55_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09234_ _18932_/Q _18931_/Q _18930_/Q vssd1 vssd1 vccd1 vccd1 _09237_/B sky130_fd_sc_hd__or3_4
XFILLER_107_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_221_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09165_ _09165_/A _10308_/A _09165_/C _09165_/D vssd1 vssd1 vccd1 vccd1 _09171_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_175_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_175_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09096_ _18800_/Q _18799_/Q _18798_/Q vssd1 vssd1 vccd1 vccd1 _09098_/C sky130_fd_sc_hd__or3_4
XFILLER_119_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_218_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_1232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09998_ _10038_/B _12066_/A vssd1 vssd1 vccd1 vccd1 _09999_/A sky130_fd_sc_hd__nor2_2
XFILLER_88_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08949_ _08967_/A vssd1 vssd1 vccd1 vccd1 _08954_/A sky130_fd_sc_hd__buf_12
XTAP_4525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_217_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11960_ _12049_/A _11960_/B _11960_/C vssd1 vssd1 vccd1 vccd1 _12028_/A sky130_fd_sc_hd__nor3_4
XFILLER_229_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10911_ _10939_/A _10443_/X _10271_/B _10903_/X _10910_/X vssd1 vssd1 vccd1 vccd1
+ _10911_/X sky130_fd_sc_hd__a41o_1
XFILLER_205_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11891_ _13418_/C vssd1 vssd1 vccd1 vccd1 _11891_/X sky130_fd_sc_hd__buf_6
XFILLER_56_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13630_ _13630_/A vssd1 vssd1 vccd1 vccd1 _13630_/X sky130_fd_sc_hd__buf_6
X_10842_ _09136_/A _09126_/B _09131_/C _09136_/C _10870_/S _10738_/A vssd1 vssd1 vccd1
+ vccd1 _10842_/X sky130_fd_sc_hd__mux4_2
XFILLER_32_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_198_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13561_ _13561_/A vssd1 vssd1 vccd1 vccd1 _13562_/A sky130_fd_sc_hd__buf_8
XFILLER_40_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10773_ _10773_/A _10773_/B _10772_/X vssd1 vssd1 vccd1 vccd1 _10773_/X sky130_fd_sc_hd__or3b_1
X_15300_ _18411_/Q _15303_/B _15299_/X _15283_/X vssd1 vssd1 vccd1 vccd1 _18411_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_40_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12512_ _11761_/A _17427_/S _12514_/A _11732_/B vssd1 vssd1 vccd1 vccd1 _12513_/B
+ sky130_fd_sc_hd__o2bb2a_1
X_16280_ _16325_/A _16285_/B vssd1 vssd1 vccd1 vccd1 _16280_/Y sky130_fd_sc_hd__nand2_1
XFILLER_200_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13492_ _13492_/A vssd1 vssd1 vccd1 vccd1 _13493_/A sky130_fd_sc_hd__buf_8
XFILLER_185_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15231_ _18432_/Q _18396_/Q _15246_/S vssd1 vssd1 vccd1 vccd1 _15231_/X sky130_fd_sc_hd__mux2_1
XFILLER_139_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12443_ _12446_/A _12493_/B vssd1 vssd1 vccd1 vccd1 _12443_/Y sky130_fd_sc_hd__nor2_1
XFILLER_60_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15162_ _15162_/A _15162_/B _15199_/C vssd1 vssd1 vccd1 vccd1 _15162_/X sky130_fd_sc_hd__or3_1
XFILLER_60_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12374_ _12381_/B _12375_/C _17894_/Q vssd1 vssd1 vccd1 vccd1 _12388_/A sky130_fd_sc_hd__o21a_1
XFILLER_165_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14113_ _12027_/A _14025_/X _14066_/X _14089_/X _14112_/X vssd1 vssd1 vccd1 vccd1
+ _14113_/X sky130_fd_sc_hd__a2111o_4
XFILLER_114_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11325_ _11323_/A _11323_/B _11339_/C vssd1 vssd1 vccd1 vccd1 _11325_/Y sky130_fd_sc_hd__o21ai_1
X_15093_ _18398_/Q _18362_/Q _15100_/S vssd1 vssd1 vccd1 vccd1 _15093_/X sky130_fd_sc_hd__mux2_1
XFILLER_154_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_180_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14044_ _18533_/Q _13857_/A _13703_/A _18548_/Q vssd1 vssd1 vccd1 vccd1 _14044_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_140_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11256_ _11922_/A _11653_/A vssd1 vssd1 vccd1 vccd1 _11257_/B sky130_fd_sc_hd__nand2_2
X_18921_ _18926_/CLK _18921_/D vssd1 vssd1 vccd1 vccd1 _18921_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_106_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10207_ _10213_/A _10213_/B _10206_/X vssd1 vssd1 vccd1 vccd1 _10217_/A sky130_fd_sc_hd__o21ai_2
XFILLER_171_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11187_ _11187_/A vssd1 vssd1 vccd1 vccd1 _17808_/D sky130_fd_sc_hd__clkbuf_1
X_18852_ _18862_/CLK _18852_/D vssd1 vssd1 vccd1 vccd1 _18852_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_79_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_228_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_171_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17803_ _17803_/CLK _17803_/D vssd1 vssd1 vccd1 vccd1 _17803_/Q sky130_fd_sc_hd__dfxtp_1
X_10138_ _18119_/Q _10138_/B vssd1 vssd1 vccd1 vccd1 _10140_/A sky130_fd_sc_hd__xnor2_2
XFILLER_171_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18783_ _18785_/CLK _18783_/D vssd1 vssd1 vccd1 vccd1 _18783_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_5760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15995_ _18612_/Q _18576_/Q _16010_/S vssd1 vssd1 vccd1 vccd1 _15995_/X sky130_fd_sc_hd__mux2_1
XFILLER_83_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17734_ _17734_/A _19012_/Q vssd1 vssd1 vccd1 vccd1 _17735_/A sky130_fd_sc_hd__and2_1
XFILLER_76_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14946_ _14949_/B _14943_/X _14945_/Y _14941_/X vssd1 vssd1 vccd1 vccd1 _18325_/D
+ sky130_fd_sc_hd__o211a_1
X_10069_ _10069_/A vssd1 vssd1 vccd1 vccd1 _10069_/X sky130_fd_sc_hd__buf_2
XFILLER_48_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_212_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17665_ _14597_/A _17663_/Y _17654_/X _17664_/Y _18978_/Q vssd1 vssd1 vccd1 vccd1
+ _17666_/B sky130_fd_sc_hd__a32o_1
XFILLER_169_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14877_ _14918_/A vssd1 vssd1 vccd1 vccd1 _14937_/B sky130_fd_sc_hd__buf_2
XINSDIODE2_101 _13848_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_112 _15162_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16616_ _16623_/B _16614_/X _16615_/X _16600_/X vssd1 vssd1 vccd1 vccd1 _18723_/D
+ sky130_fd_sc_hd__o211a_1
XINSDIODE2_123 _15233_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13828_ _12019_/A _13797_/X _13812_/X _13827_/X vssd1 vssd1 vccd1 vccd1 _13829_/D
+ sky130_fd_sc_hd__a211o_1
XFILLER_223_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINSDIODE2_134 _17120_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17596_ _17567_/X _17590_/Y _17582_/X _17592_/Y _18961_/Q vssd1 vssd1 vccd1 vccd1
+ _17597_/B sky130_fd_sc_hd__a32o_1
XFILLER_211_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_145 _15736_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_189_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_156 _18398_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_182_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16547_ _16572_/A _16551_/B vssd1 vssd1 vccd1 vccd1 _16547_/Y sky130_fd_sc_hd__nand2_1
XINSDIODE2_167 _18324_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13759_ _13759_/A vssd1 vssd1 vccd1 vccd1 _13759_/X sky130_fd_sc_hd__buf_4
XINSDIODE2_178 _17449_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_189 _09109_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_1366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16478_ _16475_/B _16474_/X _16475_/Y _16477_/X vssd1 vssd1 vccd1 vccd1 _18689_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_143_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18217_ _18217_/CLK _18217_/D vssd1 vssd1 vccd1 vccd1 _18217_/Q sky130_fd_sc_hd__dfxtp_1
X_15429_ _15431_/B _15425_/X _15426_/Y _15428_/X vssd1 vssd1 vccd1 vccd1 _18439_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_191_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19197_ _19197_/A _08982_/Y vssd1 vssd1 vccd1 vccd1 io_out[35] sky130_fd_sc_hd__ebufn_8
XFILLER_157_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18148_ _18149_/CLK _18148_/D vssd1 vssd1 vccd1 vccd1 _18148_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_145_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18079_ _18085_/CLK _18079_/D vssd1 vssd1 vccd1 vccd1 _18079_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_102_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09921_ _10278_/A vssd1 vssd1 vccd1 vccd1 _09921_/X sky130_fd_sc_hd__buf_2
XFILLER_131_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09852_ _09853_/A _09853_/B vssd1 vssd1 vccd1 vccd1 _09866_/B sky130_fd_sc_hd__xnor2_2
XTAP_541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_1307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_219_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09783_ _18111_/Q vssd1 vssd1 vccd1 vccd1 _09805_/A sky130_fd_sc_hd__clkinv_2
XTAP_596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_230_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_227_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_167_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_195_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09217_ _18674_/Q _18673_/Q _18672_/Q vssd1 vssd1 vccd1 vccd1 _09219_/C sky130_fd_sc_hd__or3_4
XFILLER_194_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_194_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09148_ _09148_/A _09148_/B _09148_/C _09148_/D vssd1 vssd1 vccd1 vccd1 _09154_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_5_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_159_1321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_147_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09079_ _09083_/A _09081_/B _17832_/Q vssd1 vssd1 vccd1 vccd1 _09080_/A sky130_fd_sc_hd__and3_1
XFILLER_194_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11110_ _11404_/A vssd1 vssd1 vccd1 vccd1 _11467_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_107_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12090_ _14247_/A _12126_/B vssd1 vssd1 vccd1 vccd1 _12095_/B sky130_fd_sc_hd__nor2_1
XFILLER_146_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11041_ _11040_/X _09742_/A _11026_/X _13370_/B vssd1 vssd1 vccd1 vccd1 _17783_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_5001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_231_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14800_ _14802_/B _14795_/X _14796_/Y _14799_/X vssd1 vssd1 vccd1 vccd1 _18289_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_5089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15780_ _15782_/B _15778_/X _15779_/Y _15763_/X vssd1 vssd1 vccd1 vccd1 _18523_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_3610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12992_ _12990_/Y _12962_/A _12951_/Y _17988_/Q _12991_/X vssd1 vssd1 vccd1 vccd1
+ _12992_/X sky130_fd_sc_hd__o221a_1
XTAP_4366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14731_ _14772_/A vssd1 vssd1 vccd1 vccd1 _14790_/B sky130_fd_sc_hd__buf_2
XFILLER_85_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_218_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11943_ _12041_/B _11947_/B _11945_/B _11945_/A _11942_/X vssd1 vssd1 vccd1 vccd1
+ _11999_/C sky130_fd_sc_hd__a221o_1
XTAP_3665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_1366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17450_ _17456_/B _17447_/X _17449_/X _17441_/X vssd1 vssd1 vccd1 vccd1 _18924_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_2942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14662_ _14687_/A _15255_/A vssd1 vssd1 vccd1 vccd1 _14670_/B sky130_fd_sc_hd__nor2_2
XTAP_3698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11874_ _11879_/A _11874_/B vssd1 vssd1 vccd1 vccd1 _17830_/D sky130_fd_sc_hd__nor2_1
XFILLER_72_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16401_ _16521_/A vssd1 vssd1 vccd1 vccd1 _16447_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_166_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13613_ _13613_/A vssd1 vssd1 vccd1 vccd1 _13738_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_77_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17381_ _17383_/B _17378_/X _17379_/Y _17380_/X vssd1 vssd1 vccd1 vccd1 _18907_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_2997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10825_ _09227_/A _09237_/B _10851_/A vssd1 vssd1 vccd1 vccd1 _10825_/X sky130_fd_sc_hd__mux2_1
XFILLER_220_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_214_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14593_ _14593_/A _17663_/A vssd1 vssd1 vccd1 vccd1 _16862_/A sky130_fd_sc_hd__or2_4
XFILLER_25_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16332_ _18690_/Q _18654_/Q _16345_/S vssd1 vssd1 vccd1 vccd1 _16332_/X sky130_fd_sc_hd__mux2_1
XFILLER_38_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13544_ _13544_/A vssd1 vssd1 vccd1 vccd1 _14016_/A sky130_fd_sc_hd__buf_4
X_10756_ _09314_/A _09319_/B _09314_/D _09314_/C _10851_/A _10856_/S vssd1 vssd1 vccd1
+ vccd1 _10757_/C sky130_fd_sc_hd__mux4_1
XFILLER_13_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_200_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16263_ _16268_/B _16259_/X _16262_/X _16252_/X vssd1 vssd1 vccd1 vccd1 _18636_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_125_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13475_ _13480_/A _13475_/B vssd1 vssd1 vccd1 vccd1 _18160_/D sky130_fd_sc_hd__nor2_1
X_10687_ _10687_/A vssd1 vssd1 vccd1 vccd1 _10695_/A sky130_fd_sc_hd__clkbuf_4
X_18002_ _18151_/CLK _18002_/D vssd1 vssd1 vccd1 vccd1 _18002_/Q sky130_fd_sc_hd__dfxtp_1
X_15214_ _15236_/A _15216_/B vssd1 vssd1 vccd1 vccd1 _15214_/Y sky130_fd_sc_hd__nand2_1
XFILLER_195_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12426_ _17900_/Q _12426_/B _12426_/C vssd1 vssd1 vccd1 vccd1 _12427_/A sky130_fd_sc_hd__and3b_1
XFILLER_103_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16194_ _16949_/A vssd1 vssd1 vccd1 vccd1 _16785_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_103_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15145_ _15145_/A _15145_/B _15145_/C vssd1 vssd1 vccd1 vccd1 _15211_/A sky130_fd_sc_hd__or3_4
XFILLER_153_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12357_ _12450_/B vssd1 vssd1 vccd1 vccd1 _12486_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_142_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11308_ _11442_/A _11655_/B _11653_/A vssd1 vssd1 vccd1 vccd1 _11308_/Y sky130_fd_sc_hd__o21ai_1
X_15076_ _15098_/A _15220_/B _15112_/C vssd1 vssd1 vccd1 vccd1 _15076_/X sky130_fd_sc_hd__or3_1
X_12288_ _12285_/C _12289_/A _11522_/A vssd1 vssd1 vccd1 vccd1 _12293_/B sky130_fd_sc_hd__o21bai_1
XFILLER_99_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14027_ _14027_/A vssd1 vssd1 vccd1 vccd1 _14027_/X sky130_fd_sc_hd__buf_6
X_18904_ _18908_/CLK _18904_/D vssd1 vssd1 vccd1 vccd1 _18904_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_214_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11239_ _11242_/B _11243_/A _11239_/C vssd1 vssd1 vccd1 vccd1 _11240_/A sky130_fd_sc_hd__and3b_1
XFILLER_45_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18835_ _18871_/CLK _18835_/D vssd1 vssd1 vccd1 vccd1 _18835_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_132_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15978_ _16000_/A _15980_/B vssd1 vssd1 vccd1 vccd1 _15978_/Y sky130_fd_sc_hd__nand2_1
X_18766_ _18773_/CLK _18766_/D vssd1 vssd1 vccd1 vccd1 _18766_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_67_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_212_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14929_ _14975_/A _15220_/B _14965_/C vssd1 vssd1 vccd1 vccd1 _14929_/X sky130_fd_sc_hd__or3_1
X_17717_ _17723_/A _19004_/Q vssd1 vssd1 vccd1 vccd1 _17718_/A sky130_fd_sc_hd__and2_1
XFILLER_110_1335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18697_ _18732_/CLK _18697_/D vssd1 vssd1 vccd1 vccd1 _18697_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_208_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_212_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17648_ _17648_/A vssd1 vssd1 vccd1 vccd1 _18974_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_1_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17579_ _17587_/A _17579_/B vssd1 vssd1 vccd1 vccd1 _17580_/A sky130_fd_sc_hd__and2_1
XFILLER_91_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_204_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_188_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_177_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09002_ _09003_/A vssd1 vssd1 vccd1 vccd1 _09002_/Y sky130_fd_sc_hd__inv_2
XFILLER_178_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_158_wb_clk_i _18114_/CLK vssd1 vssd1 vccd1 vccd1 _17990_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_105_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_172_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_160_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09904_ _09947_/A vssd1 vssd1 vccd1 vccd1 _09905_/A sky130_fd_sc_hd__buf_4
XFILLER_63_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09835_ _18100_/Q _17974_/Q vssd1 vssd1 vccd1 vccd1 _10193_/B sky130_fd_sc_hd__xor2_4
XFILLER_112_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09766_ _09816_/A _09816_/B _09816_/C vssd1 vssd1 vccd1 vccd1 _09810_/B sky130_fd_sc_hd__nand3_1
XFILLER_100_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_230_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_189_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_227_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09697_ _18263_/Q _18262_/Q _18261_/Q vssd1 vssd1 vccd1 vccd1 _09697_/X sky130_fd_sc_hd__or3_4
XFILLER_26_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_168_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_211_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10610_ _18129_/Q _10611_/B vssd1 vssd1 vccd1 vccd1 _10612_/A sky130_fd_sc_hd__and2_1
XFILLER_167_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11590_ _11984_/C _11590_/B _12023_/A vssd1 vssd1 vccd1 vccd1 _11591_/B sky130_fd_sc_hd__and3_2
XFILLER_195_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10541_ _10539_/X _10540_/X _10549_/A vssd1 vssd1 vccd1 vccd1 _10541_/X sky130_fd_sc_hd__mux2_2
XFILLER_128_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13260_ _13266_/A _18084_/Q vssd1 vssd1 vccd1 vccd1 _13261_/A sky130_fd_sc_hd__and2_1
XFILLER_210_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10472_ _10512_/B _10472_/B vssd1 vssd1 vccd1 vccd1 _10472_/X sky130_fd_sc_hd__and2_1
XFILLER_202_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12211_ _12233_/C vssd1 vssd1 vccd1 vccd1 _12239_/C sky130_fd_sc_hd__clkbuf_2
X_13191_ _13197_/A _18053_/Q vssd1 vssd1 vccd1 vccd1 _13192_/A sky130_fd_sc_hd__and2_1
XFILLER_108_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_191_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_123_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12142_ _12142_/A vssd1 vssd1 vccd1 vccd1 _13458_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_155_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16950_ _17015_/A _17528_/B _16963_/C vssd1 vssd1 vccd1 vccd1 _16950_/X sky130_fd_sc_hd__or3_1
XFILLER_123_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12073_ _12078_/A _09668_/B _12072_/X vssd1 vssd1 vccd1 vccd1 _12083_/A sky130_fd_sc_hd__a21o_1
XFILLER_46_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15901_ _15925_/A vssd1 vssd1 vccd1 vccd1 _15901_/X sky130_fd_sc_hd__clkbuf_2
X_11024_ _17971_/Q vssd1 vssd1 vccd1 vccd1 _11025_/B sky130_fd_sc_hd__buf_2
X_16881_ _18786_/Q _16884_/B _16880_/X _16871_/X vssd1 vssd1 vccd1 vccd1 _18786_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_89_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15832_ _18573_/Q _18537_/Q _15838_/S vssd1 vssd1 vccd1 vccd1 _15832_/X sky130_fd_sc_hd__mux2_1
X_18620_ _18620_/CLK _18620_/D vssd1 vssd1 vccd1 vccd1 _18620_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_66_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15763_ _15823_/A vssd1 vssd1 vccd1 vccd1 _15763_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_18551_ _18553_/CLK _18551_/D vssd1 vssd1 vccd1 vccd1 _18551_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12975_ _12975_/A _12983_/A vssd1 vssd1 vccd1 vccd1 _12976_/B sky130_fd_sc_hd__xnor2_1
XFILLER_45_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_4_2_0_wb_clk_i clkbuf_4_3_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_5_5_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_2
XTAP_3462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14714_ _18268_/Q _14715_/B _14713_/Y _14692_/X vssd1 vssd1 vccd1 vccd1 _18268_/D
+ sky130_fd_sc_hd__o211a_1
X_17502_ _17501_/B _17500_/X _17501_/Y _17497_/X vssd1 vssd1 vccd1 vccd1 _18938_/D
+ sky130_fd_sc_hd__o211a_1
X_18482_ _18482_/CLK _18482_/D vssd1 vssd1 vccd1 vccd1 _18482_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_3484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11926_ _17793_/Q _11926_/B _11951_/B vssd1 vssd1 vccd1 vccd1 _11945_/A sky130_fd_sc_hd__or3_1
X_15694_ _15694_/A _15694_/B vssd1 vssd1 vccd1 vccd1 _15694_/Y sky130_fd_sc_hd__nand2_1
XTAP_2750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_221_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17433_ _17432_/B _17431_/X _17432_/Y _17421_/X vssd1 vssd1 vccd1 vccd1 _18920_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_2772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14645_ _18253_/Q _14646_/B _14644_/Y _14629_/X vssd1 vssd1 vccd1 vccd1 _18253_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_60_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11857_ _11856_/B _11856_/C _11856_/A vssd1 vssd1 vccd1 vccd1 _11857_/Y sky130_fd_sc_hd__o21ai_1
XTAP_2794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17364_ _18939_/Q _18903_/Q _17367_/S vssd1 vssd1 vccd1 vccd1 _17364_/X sky130_fd_sc_hd__mux2_1
X_10808_ _09260_/A _09270_/D _10810_/S vssd1 vssd1 vccd1 vccd1 _10809_/B sky130_fd_sc_hd__mux2_1
X_14576_ _14598_/A vssd1 vssd1 vccd1 vccd1 _14651_/A sky130_fd_sc_hd__buf_2
XFILLER_60_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_202_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11788_ _11788_/A _11788_/B vssd1 vssd1 vccd1 vccd1 _11789_/A sky130_fd_sc_hd__nand2_1
XFILLER_158_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16315_ _16317_/B _16312_/X _16313_/Y _16314_/X vssd1 vssd1 vccd1 vccd1 _18649_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_14_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_201_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13527_ _13547_/B _13557_/A vssd1 vssd1 vccd1 vccd1 _13670_/A sky130_fd_sc_hd__nor2_4
XFILLER_159_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_203_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10739_ _10859_/S _10736_/X _10738_/X _10833_/B vssd1 vssd1 vccd1 vccd1 _10739_/X
+ sky130_fd_sc_hd__o211a_1
X_17295_ _18921_/Q _18885_/Q _17298_/S vssd1 vssd1 vccd1 vccd1 _17295_/X sky130_fd_sc_hd__mux2_1
XFILLER_9_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_220_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19034_ _19034_/CLK _19034_/D vssd1 vssd1 vccd1 vccd1 _19034_/Q sky130_fd_sc_hd__dfxtp_1
X_16246_ _16689_/A _16307_/B vssd1 vssd1 vccd1 vccd1 _16256_/B sky130_fd_sc_hd__nor2_2
XFILLER_185_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13458_ _13458_/A _13458_/B vssd1 vssd1 vccd1 vccd1 _13465_/A sky130_fd_sc_hd__or2_1
XFILLER_174_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12409_ _18990_/Q _12409_/B vssd1 vssd1 vccd1 vccd1 _12411_/B sky130_fd_sc_hd__xnor2_1
X_16177_ _16932_/A vssd1 vssd1 vccd1 vccd1 _16771_/A sky130_fd_sc_hd__buf_6
XFILLER_12_1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13389_ _13389_/A _13389_/B vssd1 vssd1 vccd1 vccd1 _13389_/Y sky130_fd_sc_hd__nand2_1
XFILLER_56_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15128_ _15178_/A _15132_/B vssd1 vssd1 vccd1 vccd1 _15128_/Y sky130_fd_sc_hd__nand2_1
XFILLER_138_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_217_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15059_ _15061_/B _15057_/X _15058_/Y _15046_/X vssd1 vssd1 vccd1 vccd1 _18352_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_68_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09620_ _18109_/Q vssd1 vssd1 vccd1 vccd1 _09645_/A sky130_fd_sc_hd__buf_2
X_18818_ _18826_/CLK _18818_/D vssd1 vssd1 vccd1 vccd1 _18818_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_68_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09551_ _09568_/A _09551_/B vssd1 vssd1 vccd1 vccd1 _09590_/B sky130_fd_sc_hd__xnor2_2
X_18749_ _18788_/CLK _18749_/D vssd1 vssd1 vccd1 vccd1 _18749_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_37_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_209_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09482_ _09482_/A _09482_/B vssd1 vssd1 vccd1 vccd1 _09483_/A sky130_fd_sc_hd__and2_1
XFILLER_23_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_197_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19118__89 vssd1 vssd1 vccd1 vccd1 _19118__89/HI _19226_/A sky130_fd_sc_hd__conb_1
XFILLER_20_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_1215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_219_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09818_ _09818_/A _09818_/B vssd1 vssd1 vccd1 vccd1 _10403_/A sky130_fd_sc_hd__xnor2_2
XFILLER_98_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_55_wb_clk_i clkbuf_5_16_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18788_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_28_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09749_ _09802_/B _09749_/B _09749_/C vssd1 vssd1 vccd1 vccd1 _09751_/A sky130_fd_sc_hd__and3_1
XFILLER_189_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_227_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_215_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12760_ _12760_/A _12947_/A _13318_/B vssd1 vssd1 vccd1 vccd1 _12760_/X sky130_fd_sc_hd__or3_1
XTAP_2035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_188_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11711_ _11619_/X _11698_/X _11707_/Y _11710_/X _11704_/C vssd1 vssd1 vccd1 vccd1
+ _11711_/X sky130_fd_sc_hd__o32a_1
XTAP_1334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12691_ _17938_/Q _12691_/B vssd1 vssd1 vccd1 vccd1 _12693_/A sky130_fd_sc_hd__xnor2_1
XFILLER_203_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_199_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14430_ _14452_/A _14430_/B vssd1 vssd1 vccd1 vccd1 _18197_/D sky130_fd_sc_hd__nor2_1
X_11642_ _17862_/Q _17861_/Q vssd1 vssd1 vccd1 vccd1 _11642_/X sky130_fd_sc_hd__or2_1
XTAP_1389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_230_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14361_ _14349_/A _14355_/C _14355_/D _14360_/X vssd1 vssd1 vccd1 vccd1 _14361_/X
+ sky130_fd_sc_hd__o31a_1
XFILLER_183_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11573_ _11573_/A vssd1 vssd1 vccd1 vccd1 _11573_/Y sky130_fd_sc_hd__inv_2
XFILLER_52_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16100_ _16701_/A _16150_/B vssd1 vssd1 vccd1 vccd1 _16109_/B sky130_fd_sc_hd__nor2_2
XFILLER_7_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13312_ _12748_/B _13318_/B _13311_/Y _12747_/B vssd1 vssd1 vccd1 vccd1 _13314_/A
+ sky130_fd_sc_hd__o31a_1
X_10524_ _09402_/A _09392_/B _09397_/C _10877_/A _10495_/S _10522_/X vssd1 vssd1 vccd1
+ vccd1 _10524_/X sky130_fd_sc_hd__mux4_1
X_17080_ _17091_/A _17080_/B vssd1 vssd1 vccd1 vccd1 _17080_/Y sky130_fd_sc_hd__nand2_1
XFILLER_182_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14292_ _14293_/A _14293_/B vssd1 vssd1 vccd1 vccd1 _14311_/A sky130_fd_sc_hd__and2_1
XFILLER_156_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16031_ _18621_/Q _18585_/Q _16031_/S vssd1 vssd1 vccd1 vccd1 _16031_/X sky130_fd_sc_hd__mux2_1
XFILLER_171_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13243_ _13243_/A vssd1 vssd1 vccd1 vccd1 _18075_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_183_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10455_ _09270_/C _09265_/D _09260_/A _09270_/D _10413_/A _10454_/X vssd1 vssd1 vccd1
+ vccd1 _10455_/X sky130_fd_sc_hd__mux4_1
XFILLER_109_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13174_ _13174_/A vssd1 vssd1 vccd1 vccd1 _18044_/D sky130_fd_sc_hd__clkbuf_1
X_10386_ _10388_/A _10386_/B vssd1 vssd1 vccd1 vccd1 _10386_/X sky130_fd_sc_hd__or2_1
XFILLER_184_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12125_ _12123_/Y _12124_/X _12099_/B _12122_/A vssd1 vssd1 vccd1 vccd1 _12127_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_97_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17982_ _17990_/CLK _17982_/D vssd1 vssd1 vccd1 vccd1 _17982_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_2_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16933_ _17514_/A _16960_/B vssd1 vssd1 vccd1 vccd1 _16943_/B sky130_fd_sc_hd__nor2_2
XFILLER_133_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12056_ _12056_/A _13649_/A vssd1 vssd1 vccd1 vccd1 _12056_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_172_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11007_ _17810_/Q vssd1 vssd1 vccd1 vccd1 _11196_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_42_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16864_ _18819_/Q _18783_/Q _16864_/S vssd1 vssd1 vccd1 vccd1 _16864_/X sky130_fd_sc_hd__mux2_1
XFILLER_203_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18603_ _18635_/CLK _18603_/D vssd1 vssd1 vccd1 vccd1 _18603_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_65_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_225_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15815_ _15815_/A _15818_/B vssd1 vssd1 vccd1 vccd1 _15815_/Y sky130_fd_sc_hd__nand2_1
XFILLER_168_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16795_ _18804_/Q _18768_/Q _16802_/S vssd1 vssd1 vccd1 vccd1 _16795_/X sky130_fd_sc_hd__mux2_1
XFILLER_206_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_206_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18534_ _18542_/CLK _18534_/D vssd1 vssd1 vccd1 vccd1 _18534_/Q sky130_fd_sc_hd__dfxtp_2
X_15746_ _18552_/Q _18516_/Q _15753_/S vssd1 vssd1 vccd1 vccd1 _15746_/X sky130_fd_sc_hd__mux2_1
XTAP_3270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12958_ _12958_/A _12958_/B vssd1 vssd1 vccd1 vccd1 _12959_/B sky130_fd_sc_hd__nor2_1
XFILLER_80_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_209_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11909_ _13526_/C vssd1 vssd1 vccd1 vccd1 _12120_/A sky130_fd_sc_hd__clkbuf_2
X_18465_ _18467_/CLK _18465_/D vssd1 vssd1 vccd1 vccd1 _18465_/Q sky130_fd_sc_hd__dfxtp_2
X_15677_ _15677_/A vssd1 vssd1 vccd1 vccd1 _15724_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_178_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12889_ _12889_/A vssd1 vssd1 vccd1 vccd1 _17959_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_209_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_221_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14628_ _14665_/A _14665_/B _15220_/B vssd1 vssd1 vccd1 vccd1 _14628_/X sky130_fd_sc_hd__or3_1
X_17416_ _18915_/Q _17419_/B _17415_/X _17400_/X vssd1 vssd1 vccd1 vccd1 _18915_/D
+ sky130_fd_sc_hd__o211a_1
X_18396_ _18398_/CLK _18396_/D vssd1 vssd1 vccd1 vccd1 _18396_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_61_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_187_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17347_ _18935_/Q _18899_/Q _17347_/S vssd1 vssd1 vccd1 vccd1 _17347_/X sky130_fd_sc_hd__mux2_1
X_14559_ _14606_/A _14559_/B vssd1 vssd1 vccd1 vccd1 _14559_/Y sky130_fd_sc_hd__nand2_1
XFILLER_119_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17278_ _18133_/Q _17278_/B vssd1 vssd1 vccd1 vccd1 _17390_/A sky130_fd_sc_hd__nand2_2
XFILLER_105_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16229_ _16268_/A _16229_/B vssd1 vssd1 vccd1 vccd1 _16229_/Y sky130_fd_sc_hd__nand2_1
X_19017_ _19019_/CLK _19017_/D vssd1 vssd1 vccd1 vccd1 _19017_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_161_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_216_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08982_ _08985_/A vssd1 vssd1 vccd1 vccd1 _08982_/Y sky130_fd_sc_hd__inv_2
XFILLER_130_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_111_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_229_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09603_ _17981_/Q vssd1 vssd1 vccd1 vccd1 _13005_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_95_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09534_ _18097_/Q _13000_/C vssd1 vssd1 vccd1 vccd1 _09535_/B sky130_fd_sc_hd__xnor2_2
XFILLER_71_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_231_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_227_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_197_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09465_ _09475_/A _09457_/B _18138_/D vssd1 vssd1 vccd1 vccd1 _18135_/D sky130_fd_sc_hd__a21o_1
XPHY_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_184_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_227_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_212_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_145_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09396_ _18365_/Q _18364_/Q _18363_/Q vssd1 vssd1 vccd1 vccd1 _09397_/D sky130_fd_sc_hd__or3_2
XFILLER_106_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_212_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_173_wb_clk_i _18114_/CLK vssd1 vssd1 vccd1 vccd1 _18088_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_149_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_1277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_102_wb_clk_i clkbuf_5_28_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18553_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_193_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_1299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_192_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_180_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10240_ _10549_/A vssd1 vssd1 vccd1 vccd1 _10923_/S sky130_fd_sc_hd__buf_4
XFILLER_191_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10171_ _10172_/A _10172_/B _10172_/C vssd1 vssd1 vccd1 vccd1 _12053_/A sky130_fd_sc_hd__a21o_1
XFILLER_79_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_1351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_219_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13930_ _18238_/Q _13544_/A _13926_/X _13929_/X vssd1 vssd1 vccd1 vccd1 _13930_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_43_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_207_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13861_ _13861_/A vssd1 vssd1 vccd1 vccd1 _13861_/X sky130_fd_sc_hd__buf_6
XFILLER_47_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15600_ _15605_/B _15598_/X _15599_/X _15595_/X vssd1 vssd1 vccd1 vccd1 _18480_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_47_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12812_ _12594_/B _17952_/Q _17957_/Q _12637_/B _12811_/X vssd1 vssd1 vccd1 vccd1
+ _12813_/D sky130_fd_sc_hd__a221o_1
X_16580_ _16780_/A vssd1 vssd1 vccd1 vccd1 _16659_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_16_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13792_ _18282_/Q _13580_/A _13734_/X _18276_/Q _13791_/X vssd1 vssd1 vccd1 vccd1
+ _13792_/X sky130_fd_sc_hd__a221o_1
XFILLER_222_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15531_ _18462_/Q _15534_/B _15530_/X _15516_/X vssd1 vssd1 vccd1 vccd1 _18462_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_103_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12743_ _12919_/B _12743_/B _12743_/C vssd1 vssd1 vccd1 vccd1 _13318_/A sky130_fd_sc_hd__and3_2
XTAP_1131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_188_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18250_ _18251_/CLK _18250_/D vssd1 vssd1 vccd1 vccd1 _18250_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_231_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15462_ _16219_/A vssd1 vssd1 vccd1 vccd1 _16055_/A sky130_fd_sc_hd__buf_4
XFILLER_163_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12674_ _17932_/Q _12635_/X _12672_/Y _12673_/X _12667_/X vssd1 vssd1 vccd1 vccd1
+ _17932_/D sky130_fd_sc_hd__a221o_1
XTAP_1186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17201_ _17200_/B _17199_/X _17200_/Y _17197_/X vssd1 vssd1 vccd1 vccd1 _18863_/D
+ sky130_fd_sc_hd__o211a_1
X_14413_ _14413_/A vssd1 vssd1 vccd1 vccd1 _18193_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_187_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11625_ _11614_/A _11339_/B _11624_/X vssd1 vssd1 vccd1 vccd1 _11625_/X sky130_fd_sc_hd__a21bo_1
X_18181_ _19000_/CLK _18181_/D vssd1 vssd1 vccd1 vccd1 _18181_/Q sky130_fd_sc_hd__dfxtp_1
X_15393_ _15993_/A _15393_/B vssd1 vssd1 vccd1 vccd1 _15403_/B sky130_fd_sc_hd__nor2_1
XFILLER_204_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17132_ _18134_/Q _17278_/B vssd1 vssd1 vccd1 vccd1 _17247_/A sky130_fd_sc_hd__nand2_2
XFILLER_11_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14344_ _14203_/X _14334_/Y _14343_/X vssd1 vssd1 vccd1 vccd1 _14344_/X sky130_fd_sc_hd__o21a_1
X_11556_ _11562_/A _12267_/A vssd1 vssd1 vccd1 vccd1 _11556_/X sky130_fd_sc_hd__or2_1
XFILLER_184_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10507_ _10559_/S vssd1 vssd1 vccd1 vccd1 _10509_/S sky130_fd_sc_hd__buf_2
X_17063_ _17068_/B _17061_/X _17062_/X _17057_/X vssd1 vssd1 vccd1 vccd1 _18828_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_171_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14275_ _14275_/A vssd1 vssd1 vccd1 vccd1 _14275_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_156_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11487_ _11784_/A _11609_/A _11453_/B _11486_/X vssd1 vssd1 vccd1 vccd1 _11488_/B
+ sky130_fd_sc_hd__o31a_1
XFILLER_183_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16014_ _16014_/A vssd1 vssd1 vccd1 vccd1 _16031_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_155_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13226_ _13226_/A vssd1 vssd1 vccd1 vccd1 _18067_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_6_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10438_ _10438_/A _14289_/A vssd1 vssd1 vccd1 vccd1 _10547_/B sky130_fd_sc_hd__nor2_2
XFILLER_139_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_100_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13157_ _13157_/A vssd1 vssd1 vccd1 vccd1 _18036_/D sky130_fd_sc_hd__clkbuf_1
XTAP_904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_174_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10369_ _09294_/A _09304_/B _10569_/A _09294_/D _10599_/S _10294_/X vssd1 vssd1 vccd1
+ vccd1 _10369_/X sky130_fd_sc_hd__mux4_1
XTAP_915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_151_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12108_ _09939_/A _09939_/B _09862_/B vssd1 vssd1 vccd1 vccd1 _12119_/A sky130_fd_sc_hd__a21o_2
XFILLER_112_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13088_ _18005_/Q _14377_/A vssd1 vssd1 vccd1 vccd1 _13089_/A sky130_fd_sc_hd__or2_1
X_17965_ _17965_/CLK _17965_/D vssd1 vssd1 vccd1 vccd1 _17965_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_112_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16916_ _16957_/A _16916_/B vssd1 vssd1 vccd1 vccd1 _16916_/Y sky130_fd_sc_hd__nand2_1
X_12039_ _12039_/A _13494_/B vssd1 vssd1 vccd1 vccd1 _12039_/X sky130_fd_sc_hd__xor2_1
XFILLER_111_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17896_ _17919_/CLK _17896_/D vssd1 vssd1 vccd1 vccd1 _17896_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_66_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16847_ _16884_/A _16847_/B vssd1 vssd1 vccd1 vccd1 _16847_/Y sky130_fd_sc_hd__nand2_1
XFILLER_92_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_225_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16778_ _18800_/Q _18764_/Q _16784_/S vssd1 vssd1 vccd1 vccd1 _16778_/X sky130_fd_sc_hd__mux2_1
XFILLER_129_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_225_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_5_11_0_wb_clk_i clkbuf_4_5_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_5_11_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_2
X_18517_ _18553_/CLK _18517_/D vssd1 vssd1 vccd1 vccd1 _18517_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_230_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15729_ _18548_/Q _18512_/Q _15733_/S vssd1 vssd1 vccd1 vccd1 _15729_/X sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_0_wb_clk_i _17929_/CLK vssd1 vssd1 vccd1 vccd1 _17954_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_222_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09250_ _18887_/Q _18886_/Q _18885_/Q vssd1 vssd1 vccd1 vccd1 _09253_/B sky130_fd_sc_hd__or3_4
XFILLER_209_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18448_ _18448_/CLK _18448_/D vssd1 vssd1 vccd1 vccd1 _18448_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_179_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_193_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09181_ _09181_/A _09181_/B _09181_/C _09181_/D vssd1 vssd1 vccd1 vccd1 _09187_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_166_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18379_ _18406_/CLK _18379_/D vssd1 vssd1 vccd1 vccd1 _18379_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_187_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_161_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_216_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08965_ _08966_/A vssd1 vssd1 vccd1 vccd1 _08965_/Y sky130_fd_sc_hd__inv_2
XFILLER_64_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_229_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_217_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09517_ _12257_/A _14383_/B _10990_/A vssd1 vssd1 vccd1 vccd1 _09517_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_227_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_212_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_197_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09448_ _09138_/B _09447_/X _09454_/B vssd1 vssd1 vccd1 vccd1 _09448_/Y sky130_fd_sc_hd__o21ai_1
XPHY_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_227_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_212_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09379_ _18380_/Q _18379_/Q _18378_/Q vssd1 vssd1 vccd1 vccd1 _09381_/C sky130_fd_sc_hd__or3_4
XFILLER_36_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11410_ _11410_/A _11546_/B vssd1 vssd1 vccd1 vccd1 _11412_/C sky130_fd_sc_hd__or2b_1
XFILLER_165_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12390_ _12390_/A vssd1 vssd1 vccd1 vccd1 _17895_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_123_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11341_ _11341_/A vssd1 vssd1 vccd1 vccd1 _11645_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_193_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_180_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14060_ _18380_/Q _13507_/A _13500_/A _18404_/Q vssd1 vssd1 vccd1 vccd1 _14060_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_125_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11272_ _11334_/A _11590_/B vssd1 vssd1 vccd1 vccd1 _11297_/B sky130_fd_sc_hd__and2_1
XFILLER_4_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13011_ _13037_/A vssd1 vssd1 vccd1 vccd1 _13011_/X sky130_fd_sc_hd__clkbuf_2
X_10223_ _10238_/A _10238_/B vssd1 vssd1 vccd1 vccd1 _10475_/A sky130_fd_sc_hd__xnor2_2
XFILLER_106_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_70_wb_clk_i clkbuf_5_20_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18696_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_3_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19102__73 vssd1 vssd1 vccd1 vccd1 _19102__73/HI _19210_/A sky130_fd_sc_hd__conb_1
XFILLER_133_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10154_ _10155_/A _13389_/A _10155_/C vssd1 vssd1 vccd1 vccd1 _10154_/X sky130_fd_sc_hd__or3_1
XTAP_5920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14962_ _14960_/B _14959_/X _14960_/Y _14961_/X vssd1 vssd1 vccd1 vccd1 _18329_/D
+ sky130_fd_sc_hd__o211a_1
X_17750_ _17756_/A _19019_/Q vssd1 vssd1 vccd1 vccd1 _17751_/A sky130_fd_sc_hd__and2_1
XFILLER_58_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10085_ _10083_/X _10084_/X _10085_/S vssd1 vssd1 vccd1 vccd1 _10086_/B sky130_fd_sc_hd__mux2_1
XTAP_5964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16701_ _16701_/A _16745_/B vssd1 vssd1 vccd1 vccd1 _16712_/B sky130_fd_sc_hd__nor2_2
XTAP_5997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13913_ _13907_/X _13912_/X _12027_/A vssd1 vssd1 vccd1 vccd1 _13913_/X sky130_fd_sc_hd__o21a_2
XFILLER_75_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14893_ _18348_/Q _18312_/Q _14905_/S vssd1 vssd1 vccd1 vccd1 _14893_/X sky130_fd_sc_hd__mux2_1
X_17681_ _17681_/A _17681_/B vssd1 vssd1 vccd1 vccd1 _17682_/A sky130_fd_sc_hd__and2_1
XFILLER_74_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_207_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_169_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16632_ _16634_/B _16630_/X _16631_/Y _16619_/X vssd1 vssd1 vccd1 vccd1 _18727_/D
+ sky130_fd_sc_hd__o211a_1
X_13844_ _18664_/Q _13539_/X _13840_/X _13843_/X vssd1 vssd1 vccd1 vccd1 _13844_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_47_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16563_ _16562_/B _16561_/X _16562_/Y _16559_/X vssd1 vssd1 vccd1 vccd1 _18710_/D
+ sky130_fd_sc_hd__o211a_1
X_13775_ _18630_/Q _13719_/X _13721_/X _18654_/Q vssd1 vssd1 vccd1 vccd1 _13775_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_16_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_222_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10987_ hold3/A _09523_/X _10977_/X _10982_/X _18995_/Q vssd1 vssd1 vccd1 vccd1 _18999_/D
+ sky130_fd_sc_hd__a32o_1
XFILLER_43_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18302_ _18307_/CLK _18302_/D vssd1 vssd1 vccd1 vccd1 _18302_/Q sky130_fd_sc_hd__dfxtp_1
X_15514_ _18495_/Q _18459_/Q _15514_/S vssd1 vssd1 vccd1 vccd1 _15514_/X sky130_fd_sc_hd__mux2_1
XFILLER_206_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12726_ _18091_/Q _18090_/Q vssd1 vssd1 vccd1 vccd1 _13322_/B sky130_fd_sc_hd__or2_1
X_16494_ _18730_/Q _18694_/Q _16509_/S vssd1 vssd1 vccd1 vccd1 _16494_/X sky130_fd_sc_hd__mux2_1
XFILLER_149_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_231_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15445_ _15445_/A _15445_/B vssd1 vssd1 vccd1 vccd1 _15445_/Y sky130_fd_sc_hd__nand2_1
X_18233_ _18809_/CLK _18233_/D vssd1 vssd1 vccd1 vccd1 _18233_/Q sky130_fd_sc_hd__dfxtp_1
X_12657_ _12656_/A _12656_/B _12591_/X vssd1 vssd1 vccd1 vccd1 _12657_/X sky130_fd_sc_hd__o21a_1
XFILLER_230_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11608_ _12233_/A _11606_/X _12235_/A _11603_/A _11615_/A vssd1 vssd1 vccd1 vccd1
+ _11608_/X sky130_fd_sc_hd__a311o_1
XFILLER_12_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15376_ _18428_/Q _15375_/B _15375_/Y _15363_/X vssd1 vssd1 vccd1 vccd1 _18428_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_157_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18164_ _18209_/CLK _18164_/D vssd1 vssd1 vccd1 vccd1 _18164_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12588_ _17925_/Q _12588_/B vssd1 vssd1 vccd1 vccd1 _12589_/A sky130_fd_sc_hd__or2_1
X_17115_ _17156_/A _17115_/B vssd1 vssd1 vccd1 vccd1 _17115_/Y sky130_fd_sc_hd__nand2_1
XFILLER_15_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14327_ _18178_/Q vssd1 vssd1 vccd1 vccd1 _16512_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_18095_ _18095_/CLK _18095_/D vssd1 vssd1 vccd1 vccd1 _18095_/Q sky130_fd_sc_hd__dfxtp_1
X_11539_ _11749_/A _11539_/B vssd1 vssd1 vccd1 vccd1 _11770_/C sky130_fd_sc_hd__nand2_2
XFILLER_8_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17046_ _17091_/A _17046_/B vssd1 vssd1 vccd1 vccd1 _17046_/Y sky130_fd_sc_hd__nand2_1
X_14258_ _14317_/A _09711_/A _10679_/X _14237_/X vssd1 vssd1 vccd1 vccd1 _14258_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_144_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_217_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13209_ _13209_/A vssd1 vssd1 vccd1 vccd1 _18060_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_87_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14189_ _14332_/S _18994_/Q _14330_/B vssd1 vssd1 vccd1 vccd1 _14355_/D sky130_fd_sc_hd__nor3_2
XTAP_712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18997_ _18997_/CLK _18997_/D vssd1 vssd1 vccd1 vccd1 _18997_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_26_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17948_ _17954_/CLK _17948_/D vssd1 vssd1 vccd1 vccd1 _17948_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_22_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_215_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_227_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_226_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17879_ _17879_/CLK _17879_/D vssd1 vssd1 vccd1 vccd1 _17879_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_227_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_226_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_226_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09302_ _18485_/Q _18484_/Q _18483_/Q vssd1 vssd1 vccd1 vccd1 _09304_/C sky130_fd_sc_hd__or3_2
XFILLER_22_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_224_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_221_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_210_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09233_ _18929_/Q _18928_/Q _18927_/Q vssd1 vssd1 vccd1 vccd1 _09237_/A sky130_fd_sc_hd__or3_4
XFILLER_22_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_4_15_0_wb_clk_i clkbuf_3_7_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_5_31_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_2
X_09164_ _18644_/Q _18643_/Q _18642_/Q vssd1 vssd1 vccd1 vccd1 _09165_/D sky130_fd_sc_hd__or3_4
XFILLER_33_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09095_ _18773_/Q _18772_/Q _18771_/Q vssd1 vssd1 vccd1 vccd1 _09098_/B sky130_fd_sc_hd__or3_4
XFILLER_119_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_123_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_142_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09997_ _10942_/A _09989_/X _09996_/X _09694_/A vssd1 vssd1 vccd1 vccd1 _09997_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_49_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08948_ _08948_/A vssd1 vssd1 vccd1 vccd1 _08948_/Y sky130_fd_sc_hd__inv_2
XTAP_4515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_229_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10910_ _14330_/A _10910_/B _10910_/C _10910_/D vssd1 vssd1 vccd1 vccd1 _10910_/X
+ sky130_fd_sc_hd__and4b_1
XTAP_3858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11890_ _12224_/A vssd1 vssd1 vccd1 vccd1 _13418_/C sky130_fd_sc_hd__buf_6
XFILLER_72_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10841_ _10841_/A vssd1 vssd1 vccd1 vccd1 _10870_/S sky130_fd_sc_hd__buf_4
XFILLER_204_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13560_ _13560_/A vssd1 vssd1 vccd1 vccd1 _13561_/A sky130_fd_sc_hd__buf_8
XFILLER_44_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10772_ _10838_/A _10818_/B _10772_/C vssd1 vssd1 vccd1 vccd1 _10772_/X sky130_fd_sc_hd__or3_1
XFILLER_213_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12511_ _12509_/A _17427_/S _12509_/Y _12510_/X vssd1 vssd1 vccd1 vccd1 _17912_/D
+ sky130_fd_sc_hd__a211o_1
XFILLER_157_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13491_ _13857_/A vssd1 vssd1 vccd1 vccd1 _13492_/A sky130_fd_sc_hd__buf_6
XFILLER_12_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15230_ _15250_/A vssd1 vssd1 vccd1 vccd1 _15246_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_185_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12442_ _17902_/Q vssd1 vssd1 vccd1 vccd1 _12446_/A sky130_fd_sc_hd__inv_2
XFILLER_12_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15161_ _18414_/Q _18378_/Q _15177_/S vssd1 vssd1 vccd1 vccd1 _15161_/X sky130_fd_sc_hd__mux2_1
XFILLER_5_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12373_ _12373_/A _18987_/Q vssd1 vssd1 vccd1 vccd1 _12375_/C sky130_fd_sc_hd__and2_1
XFILLER_125_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14112_ _12028_/D _14096_/X _14111_/X vssd1 vssd1 vccd1 vccd1 _14112_/X sky130_fd_sc_hd__a21o_1
XFILLER_125_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11324_ _17878_/Q _19030_/Q vssd1 vssd1 vccd1 vccd1 _11339_/C sky130_fd_sc_hd__nor2b_2
XFILLER_5_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15092_ _15094_/B _15090_/X _15091_/Y _15083_/X vssd1 vssd1 vccd1 vccd1 _18361_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_158_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_181_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14043_ _18551_/Q _13838_/A _14017_/A _18527_/Q vssd1 vssd1 vccd1 vccd1 _14043_/X
+ sky130_fd_sc_hd__a22o_1
X_18920_ _18959_/CLK _18920_/D vssd1 vssd1 vccd1 vccd1 _18920_/Q sky130_fd_sc_hd__dfxtp_4
X_11255_ _11735_/B vssd1 vssd1 vccd1 vccd1 _11748_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_106_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10206_ _10206_/A _10206_/B vssd1 vssd1 vccd1 vccd1 _10206_/X sky130_fd_sc_hd__or2_1
X_18851_ _18865_/CLK _18851_/D vssd1 vssd1 vccd1 vccd1 _18851_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_136_1355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11186_ _11196_/D _11198_/B _11186_/C vssd1 vssd1 vccd1 vccd1 _11187_/A sky130_fd_sc_hd__and3b_1
XFILLER_192_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17802_ _17851_/CLK _17802_/D vssd1 vssd1 vccd1 vccd1 _17802_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_79_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_171_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10137_ _10135_/X _10137_/B vssd1 vssd1 vccd1 vccd1 _10138_/B sky130_fd_sc_hd__and2b_1
XFILLER_95_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18782_ _18821_/CLK _18782_/D vssd1 vssd1 vccd1 vccd1 _18782_/Q sky130_fd_sc_hd__dfxtp_4
XTAP_5750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15994_ _16014_/A vssd1 vssd1 vccd1 vccd1 _16010_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_121_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17733_ _17733_/A vssd1 vssd1 vccd1 vccd1 _19010_/D sky130_fd_sc_hd__clkbuf_1
X_14945_ _14992_/A _14949_/B vssd1 vssd1 vccd1 vccd1 _14945_/Y sky130_fd_sc_hd__nand2_1
X_10068_ _12063_/A _14317_/B _10068_/C vssd1 vssd1 vccd1 vccd1 _10068_/X sky130_fd_sc_hd__and3_1
XTAP_5794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_205_wb_clk_i clkbuf_5_6_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18977_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_76_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17664_ _17663_/Y _17604_/X _14386_/A vssd1 vssd1 vccd1 vccd1 _17664_/Y sky130_fd_sc_hd__a21oi_1
X_14876_ _14875_/B _14874_/X _14875_/Y _14859_/X vssd1 vssd1 vccd1 vccd1 _18308_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_211_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINSDIODE2_102 _13858_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_169_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16615_ _16615_/A _16759_/B _16628_/C vssd1 vssd1 vccd1 vccd1 _16615_/X sky130_fd_sc_hd__or3_1
XINSDIODE2_113 _15162_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XINSDIODE2_124 _15243_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13827_ _12027_/D _13819_/X _13826_/X _12022_/C vssd1 vssd1 vccd1 vccd1 _13827_/X
+ sky130_fd_sc_hd__a22o_1
X_17595_ _17595_/A vssd1 vssd1 vccd1 vccd1 _18960_/D sky130_fd_sc_hd__clkbuf_1
XINSDIODE2_135 _17120_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_204_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_146 _16749_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_189_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_157 _18342_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16546_ _18742_/Q _18706_/Q _16546_/S vssd1 vssd1 vccd1 vccd1 _16546_/X sky130_fd_sc_hd__mux2_1
X_13758_ _13758_/A vssd1 vssd1 vccd1 vccd1 _13759_/A sky130_fd_sc_hd__buf_6
XINSDIODE2_168 _18329_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_210_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_179 _17736_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_206_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_203_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_189_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12709_ _12709_/A vssd1 vssd1 vccd1 vccd1 _17937_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_91_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16477_ _16559_/A vssd1 vssd1 vccd1 vccd1 _16477_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_13689_ _18594_/Q _13505_/A _13626_/A _18618_/Q vssd1 vssd1 vccd1 vccd1 _13689_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_86_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18216_ _18217_/CLK _18216_/D vssd1 vssd1 vccd1 vccd1 _18216_/Q sky130_fd_sc_hd__dfxtp_1
X_15428_ _15516_/A vssd1 vssd1 vccd1 vccd1 _15428_/X sky130_fd_sc_hd__clkbuf_2
X_19196_ _19196_/A _08981_/Y vssd1 vssd1 vccd1 vccd1 io_out[34] sky130_fd_sc_hd__ebufn_8
XFILLER_54_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15359_ _15366_/B _15356_/X _15358_/X _15340_/X vssd1 vssd1 vccd1 vccd1 _18423_/D
+ sky130_fd_sc_hd__o211a_1
X_18147_ _18147_/CLK _18147_/D vssd1 vssd1 vccd1 vccd1 _18147_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_157_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18078_ _18085_/CLK _18078_/D vssd1 vssd1 vccd1 vccd1 _18078_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_105_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09920_ _12122_/A _09920_/B vssd1 vssd1 vccd1 vccd1 _10278_/A sky130_fd_sc_hd__and2_2
XFILLER_160_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17029_ _17035_/B _17026_/X _17028_/X _17020_/X vssd1 vssd1 vccd1 vccd1 _18819_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_144_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_1305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09851_ _18101_/Q _10627_/B _09850_/X vssd1 vssd1 vccd1 vccd1 _09853_/B sky130_fd_sc_hd__a21oi_2
XFILLER_112_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_213_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09782_ _17784_/Q _09779_/X _09780_/Y _09781_/Y vssd1 vssd1 vccd1 vccd1 _09891_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_100_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_218_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19093__64 vssd1 vssd1 vccd1 vccd1 _19093__64/HI _19201_/A sky130_fd_sc_hd__conb_1
XTAP_586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_227_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_227_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_227_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_226_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_228_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_224_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09216_ _18686_/Q _18685_/Q _18684_/Q vssd1 vssd1 vccd1 vccd1 _09219_/B sky130_fd_sc_hd__or3_4
XFILLER_10_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09147_ _18725_/Q _18724_/Q _18723_/Q vssd1 vssd1 vccd1 vccd1 _09148_/D sky130_fd_sc_hd__or3_4
XFILLER_33_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_5_4_0_wb_clk_i clkbuf_5_5_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_5_4_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_68_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09078_ _09078_/A vssd1 vssd1 vccd1 vccd1 _19185_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_159_1366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11040_ _13344_/A vssd1 vssd1 vccd1 vccd1 _11040_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_89_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12991_ _12760_/A _13019_/B _13318_/C _12927_/Y vssd1 vssd1 vccd1 vccd1 _12991_/X
+ sky130_fd_sc_hd__o31a_2
XFILLER_40_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14730_ _14729_/B _14728_/X _14729_/Y _14716_/X vssd1 vssd1 vccd1 vccd1 _18272_/D
+ sky130_fd_sc_hd__o211a_1
X_11942_ _11942_/A _17787_/Q _17786_/Q _17785_/Q vssd1 vssd1 vccd1 vccd1 _11942_/X
+ sky130_fd_sc_hd__or4_2
XFILLER_229_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_1326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14661_ _16932_/A vssd1 vssd1 vccd1 vccd1 _15255_/A sky130_fd_sc_hd__buf_6
XTAP_3688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11873_ hold1/X _11867_/X _11870_/Y vssd1 vssd1 vccd1 vccd1 _11874_/B sky130_fd_sc_hd__a21oi_1
XTAP_2954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16400_ _18706_/Q _18670_/Q _16400_/S vssd1 vssd1 vccd1 vccd1 _16400_/X sky130_fd_sc_hd__mux2_1
X_13612_ _13612_/A vssd1 vssd1 vccd1 vccd1 _13612_/X sky130_fd_sc_hd__buf_6
XFILLER_38_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10824_ _10824_/A vssd1 vssd1 vccd1 vccd1 _12092_/A sky130_fd_sc_hd__buf_4
XFILLER_60_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14592_ _14609_/B vssd1 vssd1 vccd1 vccd1 _17663_/A sky130_fd_sc_hd__clkbuf_2
X_17380_ _17400_/A vssd1 vssd1 vccd1 vccd1 _17380_/X sky130_fd_sc_hd__clkbuf_2
XTAP_2998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_207_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16331_ _16771_/A _16356_/B vssd1 vssd1 vccd1 vccd1 _16342_/B sky130_fd_sc_hd__nor2_2
XFILLER_186_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13543_ _13749_/A vssd1 vssd1 vccd1 vccd1 _13544_/A sky130_fd_sc_hd__clkbuf_4
X_10755_ _10877_/B vssd1 vssd1 vccd1 vccd1 _10851_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_38_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16262_ _16310_/A _16703_/B _16272_/C vssd1 vssd1 vccd1 vccd1 _16262_/X sky130_fd_sc_hd__or3_1
XFILLER_186_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13474_ _17844_/Q _13464_/X _13465_/X vssd1 vssd1 vccd1 vccd1 _13475_/B sky130_fd_sc_hd__a21oi_1
XFILLER_186_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10686_ _10716_/A vssd1 vssd1 vccd1 vccd1 _10687_/A sky130_fd_sc_hd__buf_6
X_15213_ _18390_/Q _15216_/B _15212_/X _15208_/X vssd1 vssd1 vccd1 vccd1 _18390_/D
+ sky130_fd_sc_hd__o211a_1
X_18001_ _18088_/CLK _18001_/D vssd1 vssd1 vccd1 vccd1 _18001_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_173_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12425_ _18991_/Q vssd1 vssd1 vccd1 vccd1 _12426_/B sky130_fd_sc_hd__inv_2
X_16193_ _16193_/A vssd1 vssd1 vccd1 vccd1 _16248_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_200_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15144_ _15142_/B _15141_/X _15142_/Y _15143_/X vssd1 vssd1 vccd1 vccd1 _18374_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_138_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12356_ _12420_/B vssd1 vssd1 vccd1 vccd1 _12450_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_181_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_181_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11307_ _11403_/A _11307_/B vssd1 vssd1 vccd1 vccd1 _11655_/B sky130_fd_sc_hd__and2_2
XFILLER_4_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15075_ _18393_/Q _18357_/Q _15081_/S vssd1 vssd1 vccd1 vccd1 _15075_/X sky130_fd_sc_hd__mux2_1
XFILLER_5_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12287_ _12287_/A _12304_/A vssd1 vssd1 vccd1 vccd1 _12287_/Y sky130_fd_sc_hd__nor2_1
XFILLER_206_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14026_ _14026_/A vssd1 vssd1 vccd1 vccd1 _14027_/A sky130_fd_sc_hd__buf_6
X_18903_ _18908_/CLK _18903_/D vssd1 vssd1 vccd1 vccd1 _18903_/Q sky130_fd_sc_hd__dfxtp_2
X_11238_ _11237_/B _11232_/C _11892_/A vssd1 vssd1 vccd1 vccd1 _11239_/C sky130_fd_sc_hd__a21o_1
XFILLER_175_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18834_ _18871_/CLK _18834_/D vssd1 vssd1 vccd1 vccd1 _18834_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_171_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11169_ _17806_/Q _11169_/B _11169_/C _17808_/Q vssd1 vssd1 vccd1 vccd1 _11169_/X
+ sky130_fd_sc_hd__or4b_1
XFILLER_67_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18765_ _18765_/CLK _18765_/D vssd1 vssd1 vccd1 vccd1 _18765_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_5580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15977_ _18570_/Q _15980_/B _15976_/X _15972_/X vssd1 vssd1 vccd1 vccd1 _18570_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_222_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_212_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17716_ _17716_/A vssd1 vssd1 vccd1 vccd1 _19002_/D sky130_fd_sc_hd__clkbuf_1
X_14928_ _14928_/A vssd1 vssd1 vccd1 vccd1 _14975_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_18696_ _18696_/CLK _18696_/D vssd1 vssd1 vccd1 vccd1 _18696_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_36_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_1347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_224_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_223_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17647_ _17659_/A _17647_/B vssd1 vssd1 vccd1 vccd1 _17648_/A sky130_fd_sc_hd__and2_1
XFILLER_224_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14859_ _14881_/A vssd1 vssd1 vccd1 vccd1 _14859_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_21_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_212_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_205_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17578_ _17575_/X _17576_/Y _17561_/X _17577_/Y _18957_/Q vssd1 vssd1 vccd1 vccd1
+ _17579_/B sky130_fd_sc_hd__a32o_1
XFILLER_50_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_149_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16529_ _16641_/A vssd1 vssd1 vccd1 vccd1 _16621_/A sky130_fd_sc_hd__buf_2
XFILLER_108_1243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09001_ _09003_/A vssd1 vssd1 vccd1 vccd1 _09001_/Y sky130_fd_sc_hd__inv_2
XFILLER_192_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19179_ _19179_/A _09012_/Y vssd1 vssd1 vccd1 vccd1 io_out[17] sky130_fd_sc_hd__ebufn_8
XFILLER_118_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_105_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_1271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09903_ _10294_/A vssd1 vssd1 vccd1 vccd1 _09947_/A sky130_fd_sc_hd__clkbuf_4
Xclkbuf_leaf_198_wb_clk_i _18176_/CLK vssd1 vssd1 vccd1 vccd1 _18184_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_28_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_127_wb_clk_i clkbuf_5_24_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18387_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_63_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09834_ _11032_/A _09834_/B vssd1 vssd1 vccd1 vccd1 _09839_/A sky130_fd_sc_hd__xnor2_4
XFILLER_24_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09765_ _09792_/A _09792_/B vssd1 vssd1 vccd1 vccd1 _09816_/C sky130_fd_sc_hd__or2_1
XFILLER_6_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_227_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_230_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09696_ _18242_/Q _18241_/Q _18240_/Q vssd1 vssd1 vccd1 vccd1 _09696_/X sky130_fd_sc_hd__or3_4
XTAP_2206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_227_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_214_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_1340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10540_ _09715_/X _09714_/X _09713_/X _09712_/X _10522_/A _10509_/S vssd1 vssd1 vccd1
+ vccd1 _10540_/X sky130_fd_sc_hd__mux4_1
XFILLER_194_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_202_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10471_ _10469_/X _10470_/X _10902_/S vssd1 vssd1 vccd1 vccd1 _10472_/B sky130_fd_sc_hd__mux2_2
XFILLER_182_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_157_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12210_ _12210_/A _12210_/B vssd1 vssd1 vccd1 vccd1 _12233_/C sky130_fd_sc_hd__or2_2
XFILLER_202_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13190_ _13190_/A vssd1 vssd1 vccd1 vccd1 _18051_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_203_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_191_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12141_ _12141_/A _12141_/B vssd1 vssd1 vccd1 vccd1 _12180_/B sky130_fd_sc_hd__nand2_1
XFILLER_11_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_194_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_150_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_172_1330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12072_ _09667_/B _12072_/B vssd1 vssd1 vccd1 vccd1 _12072_/X sky130_fd_sc_hd__and2b_1
XFILLER_96_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15900_ _15942_/A _15900_/B vssd1 vssd1 vccd1 vccd1 _15900_/Y sky130_fd_sc_hd__nand2_1
XFILLER_2_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11023_ _11023_/A vssd1 vssd1 vccd1 vccd1 _11023_/X sky130_fd_sc_hd__buf_4
XFILLER_42_1208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16880_ _16936_/A _16880_/B _16936_/C vssd1 vssd1 vccd1 vccd1 _16880_/X sky130_fd_sc_hd__or3_1
XFILLER_2_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15831_ _15982_/A _15844_/B vssd1 vssd1 vccd1 vccd1 _15839_/B sky130_fd_sc_hd__nor2_1
XTAP_4120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18550_ _18553_/CLK _18550_/D vssd1 vssd1 vccd1 vccd1 _18550_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15762_ _15799_/A _15909_/B _15811_/C vssd1 vssd1 vccd1 vccd1 _15762_/X sky130_fd_sc_hd__or3_1
XTAP_4175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12974_ _12967_/A _12958_/B _12970_/A vssd1 vssd1 vccd1 vccd1 _12976_/A sky130_fd_sc_hd__a21o_1
XFILLER_206_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17501_ _17512_/A _17501_/B vssd1 vssd1 vccd1 vccd1 _17501_/Y sky130_fd_sc_hd__nand2_1
XTAP_3463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14713_ _14750_/A _14715_/B vssd1 vssd1 vccd1 vccd1 _14713_/Y sky130_fd_sc_hd__nand2_1
XFILLER_46_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18481_ _18482_/CLK _18481_/D vssd1 vssd1 vccd1 vccd1 _18481_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11925_ _11925_/A _12126_/B vssd1 vssd1 vccd1 vccd1 _11925_/X sky130_fd_sc_hd__or2_1
X_15693_ _18539_/Q _18503_/Q _15693_/S vssd1 vssd1 vccd1 vccd1 _15693_/X sky130_fd_sc_hd__mux2_1
XFILLER_206_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17432_ _17456_/A _17432_/B vssd1 vssd1 vccd1 vccd1 _17432_/Y sky130_fd_sc_hd__nand2_1
XTAP_2773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14644_ _14681_/A _14646_/B vssd1 vssd1 vccd1 vccd1 _14644_/Y sky130_fd_sc_hd__nand2_1
X_11856_ _11856_/A _11856_/B _11856_/C vssd1 vssd1 vccd1 vccd1 _11856_/X sky130_fd_sc_hd__or3_1
XFILLER_162_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_214_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10807_ _10798_/X _10802_/X _10806_/X _10707_/Y vssd1 vssd1 vccd1 vccd1 _10822_/B
+ sky130_fd_sc_hd__o211a_1
X_14575_ _18239_/Q _14574_/B _14574_/Y _14561_/X vssd1 vssd1 vccd1 vccd1 _18239_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_20_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17363_ _17503_/A _17397_/B vssd1 vssd1 vccd1 vccd1 _17372_/B sky130_fd_sc_hd__nor2_2
X_11787_ _11542_/B _11788_/B _11795_/B vssd1 vssd1 vccd1 vccd1 _11787_/X sky130_fd_sc_hd__o21a_1
XFILLER_13_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16314_ _16354_/A vssd1 vssd1 vccd1 vccd1 _16314_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_202_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10738_ _10738_/A _10738_/B vssd1 vssd1 vccd1 vccd1 _10738_/X sky130_fd_sc_hd__or2_1
XFILLER_9_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13526_ _13526_/A _13526_/B _13526_/C vssd1 vssd1 vccd1 vccd1 _13547_/B sky130_fd_sc_hd__or3_4
XFILLER_201_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17294_ _17435_/A _17351_/B vssd1 vssd1 vccd1 vccd1 _17303_/B sky130_fd_sc_hd__nor2_2
XFILLER_146_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19033_ _19035_/CLK _19033_/D vssd1 vssd1 vccd1 vccd1 _19033_/Q sky130_fd_sc_hd__dfxtp_1
X_16245_ _16289_/A vssd1 vssd1 vccd1 vccd1 _16307_/B sky130_fd_sc_hd__buf_2
X_13457_ _13457_/A vssd1 vssd1 vccd1 vccd1 _13457_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_220_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10669_ _10737_/S vssd1 vssd1 vccd1 vccd1 _10882_/S sky130_fd_sc_hd__buf_4
XFILLER_12_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12408_ _12408_/A vssd1 vssd1 vccd1 vccd1 _17897_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_51_1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16176_ _16175_/B _16174_/X _16175_/Y _16162_/X vssd1 vssd1 vccd1 vccd1 _18617_/D
+ sky130_fd_sc_hd__o211a_1
X_13388_ _18118_/Q _13344_/X _13342_/X _13383_/X vssd1 vssd1 vccd1 vccd1 _18118_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_142_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15127_ _15247_/A vssd1 vssd1 vccd1 vccd1 _15178_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_126_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12339_ _17888_/Q _11463_/B _12336_/X vssd1 vssd1 vccd1 vccd1 _12340_/C sky130_fd_sc_hd__a21oi_2
XFILLER_99_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_217_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15058_ _15058_/A _15061_/B vssd1 vssd1 vccd1 vccd1 _15058_/Y sky130_fd_sc_hd__nand2_1
XFILLER_99_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14009_ _14009_/A _14009_/B _14009_/C _14009_/D vssd1 vssd1 vccd1 vccd1 _14009_/X
+ sky130_fd_sc_hd__or4_1
XFILLER_96_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_214_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18817_ _18826_/CLK _18817_/D vssd1 vssd1 vccd1 vccd1 _18817_/Q sky130_fd_sc_hd__dfxtp_2
X_19063__34 vssd1 vssd1 vccd1 vccd1 _19063__34/HI _19157_/A sky130_fd_sc_hd__conb_1
XFILLER_3_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09550_ _10142_/A _09570_/B vssd1 vssd1 vccd1 vccd1 _09551_/B sky130_fd_sc_hd__xor2_1
X_18748_ _18752_/CLK _18748_/D vssd1 vssd1 vccd1 vccd1 _18748_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_3_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09481_ _09463_/X _09482_/B _18146_/D vssd1 vssd1 vccd1 vccd1 _18147_/D sky130_fd_sc_hd__o21a_1
X_18679_ _18682_/CLK _18679_/D vssd1 vssd1 vccd1 vccd1 _18679_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_52_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_224_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_225_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_165_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_1262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_1355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_219_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_219_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09817_ _09817_/A _09817_/B vssd1 vssd1 vccd1 vccd1 _09818_/B sky130_fd_sc_hd__nor2_1
XFILLER_74_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09748_ _09748_/A _09753_/A _09748_/C vssd1 vssd1 vccd1 vccd1 _09749_/C sky130_fd_sc_hd__nand3_1
XFILLER_185_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_1274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09679_ _09679_/A _09649_/X vssd1 vssd1 vccd1 vccd1 _09699_/B sky130_fd_sc_hd__nor2b_4
XFILLER_28_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_95_wb_clk_i _18254_/CLK vssd1 vssd1 vccd1 vccd1 _18251_/CLK sky130_fd_sc_hd__clkbuf_16
X_11710_ _11390_/X _11698_/X _11708_/Y _11709_/X _11619_/X vssd1 vssd1 vccd1 vccd1
+ _11710_/X sky130_fd_sc_hd__o32a_1
XFILLER_42_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12690_ _17934_/Q _12613_/A _12688_/Y _12689_/X _12667_/X vssd1 vssd1 vccd1 vccd1
+ _17934_/D sky130_fd_sc_hd__a221o_1
XFILLER_153_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_24_wb_clk_i clkbuf_5_6_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18959_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_11641_ _17863_/Q _19035_/Q vssd1 vssd1 vccd1 vccd1 _11651_/A sky130_fd_sc_hd__and2b_1
XFILLER_42_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14360_ _18184_/Q vssd1 vssd1 vccd1 vccd1 _14360_/X sky130_fd_sc_hd__buf_4
X_11572_ _12261_/A _11390_/A _11566_/Y _11571_/Y _11619_/A vssd1 vssd1 vccd1 vccd1
+ _11573_/A sky130_fd_sc_hd__o32a_1
XFILLER_211_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_183_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13311_ _13311_/A _13311_/B _13311_/C _13311_/D vssd1 vssd1 vccd1 vccd1 _13311_/Y
+ sky130_fd_sc_hd__nor4_2
X_10523_ _09402_/D _09397_/D _09392_/C _09397_/B _10495_/S _10522_/X vssd1 vssd1 vccd1
+ vccd1 _10523_/X sky130_fd_sc_hd__mux4_1
XFILLER_122_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_196_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_183_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14291_ _14319_/S _12130_/A _14289_/Y _14290_/X vssd1 vssd1 vccd1 vccd1 _14293_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_202_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16030_ _16030_/A _16041_/B vssd1 vssd1 vccd1 vccd1 _16039_/B sky130_fd_sc_hd__nor2_2
X_13242_ _13244_/A _18076_/Q vssd1 vssd1 vccd1 vccd1 _13243_/A sky130_fd_sc_hd__and2_1
XFILLER_108_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10454_ _10498_/A vssd1 vssd1 vccd1 vccd1 _10454_/X sky130_fd_sc_hd__buf_4
XFILLER_6_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13173_ _13175_/A _18045_/Q vssd1 vssd1 vccd1 vccd1 _13174_/A sky130_fd_sc_hd__and2_1
XFILLER_184_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10385_ _09314_/B _09319_/A _09319_/C _09309_/C _09972_/B _09905_/A vssd1 vssd1 vccd1
+ vccd1 _10386_/B sky130_fd_sc_hd__mux4_2
XFILLER_123_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12124_ _12124_/A _13526_/A vssd1 vssd1 vccd1 vccd1 _12124_/X sky130_fd_sc_hd__or2_1
XFILLER_184_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17981_ _17990_/CLK _17981_/D vssd1 vssd1 vccd1 vccd1 _17981_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_2_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16932_ _16932_/A vssd1 vssd1 vccd1 vccd1 _17514_/A sky130_fd_sc_hd__buf_6
X_12055_ _12055_/A _12055_/B _12055_/C _12055_/D vssd1 vssd1 vccd1 vccd1 _13649_/A
+ sky130_fd_sc_hd__nor4_4
XFILLER_46_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11006_ _17812_/Q vssd1 vssd1 vccd1 vccd1 _11201_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_38_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16863_ _17458_/A _16906_/B vssd1 vssd1 vccd1 vccd1 _16874_/B sky130_fd_sc_hd__nor2_2
XFILLER_226_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18602_ _18608_/CLK _18602_/D vssd1 vssd1 vccd1 vccd1 _18602_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_65_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15814_ _18568_/Q _18532_/Q _15838_/S vssd1 vssd1 vccd1 vccd1 _15814_/X sky130_fd_sc_hd__mux2_1
XFILLER_219_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16794_ _16794_/A _16794_/B vssd1 vssd1 vccd1 vccd1 _16803_/B sky130_fd_sc_hd__nor2_2
XFILLER_65_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_225_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18533_ _18533_/CLK _18533_/D vssd1 vssd1 vccd1 vccd1 _18533_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_19_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15745_ _16041_/A _15745_/B vssd1 vssd1 vccd1 vccd1 _15754_/B sky130_fd_sc_hd__nor2_1
XTAP_3260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12957_ _12958_/A _12958_/B vssd1 vssd1 vccd1 vccd1 _12969_/A sky130_fd_sc_hd__and2_1
XFILLER_45_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18464_ _18485_/CLK _18464_/D vssd1 vssd1 vccd1 vccd1 _18464_/Q sky130_fd_sc_hd__dfxtp_1
X_11908_ _17804_/Q _12037_/A vssd1 vssd1 vccd1 vccd1 _13526_/C sky130_fd_sc_hd__xnor2_4
X_15676_ _16287_/A _15748_/C vssd1 vssd1 vccd1 vccd1 _15683_/B sky130_fd_sc_hd__nor2_1
XFILLER_206_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12888_ _12890_/B _12888_/B _12888_/C vssd1 vssd1 vccd1 vccd1 _12889_/A sky130_fd_sc_hd__and3b_1
XTAP_2581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17415_ _17437_/A _17415_/B _17460_/C vssd1 vssd1 vccd1 vccd1 _17415_/X sky130_fd_sc_hd__or3_1
X_14627_ _16889_/A vssd1 vssd1 vccd1 vccd1 _15220_/B sky130_fd_sc_hd__buf_6
X_18395_ _18398_/CLK _18395_/D vssd1 vssd1 vccd1 vccd1 _18395_/Q sky130_fd_sc_hd__dfxtp_2
X_11839_ _11491_/A _11371_/B _11833_/X _11838_/X _11501_/X vssd1 vssd1 vccd1 vccd1
+ _11842_/B sky130_fd_sc_hd__o311a_1
XTAP_1880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17346_ _17349_/B _17343_/X _17345_/Y _17341_/X vssd1 vssd1 vccd1 vccd1 _18898_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_158_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14558_ _18235_/Q _14559_/B _14557_/Y _14533_/X vssd1 vssd1 vccd1 vccd1 _18235_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_14_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13509_ _13509_/A _13509_/B vssd1 vssd1 vccd1 vccd1 _13563_/A sky130_fd_sc_hd__nand2_8
XFILLER_173_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_1208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17277_ _17423_/A _17399_/C vssd1 vssd1 vccd1 vccd1 _17291_/B sky130_fd_sc_hd__nor2_2
XFILLER_174_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14489_ _18219_/Q _14491_/B vssd1 vssd1 vccd1 vccd1 _14490_/A sky130_fd_sc_hd__and2_1
XFILLER_220_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19016_ _19029_/CLK _19016_/D vssd1 vssd1 vccd1 vccd1 _19016_/Q sky130_fd_sc_hd__dfxtp_1
X_16228_ _18628_/Q _16229_/B _16227_/Y _16209_/X vssd1 vssd1 vccd1 vccd1 _18628_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_174_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16159_ _18650_/Q _18614_/Q _16170_/S vssd1 vssd1 vccd1 vccd1 _16159_/X sky130_fd_sc_hd__mux2_1
XFILLER_127_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08981_ _08985_/A vssd1 vssd1 vccd1 vccd1 _08981_/Y sky130_fd_sc_hd__inv_2
XFILLER_130_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_218_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_1293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09602_ _10123_/A vssd1 vssd1 vccd1 vccd1 _10124_/A sky130_fd_sc_hd__inv_2
XFILLER_216_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09533_ _17978_/Q vssd1 vssd1 vccd1 vccd1 _13000_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_3_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_184_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09464_ _09463_/X _09461_/A _18134_/D vssd1 vssd1 vccd1 vccd1 _18133_/D sky130_fd_sc_hd__a21o_1
XFILLER_36_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_227_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_184_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_212_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09395_ _18344_/Q _18343_/Q _18342_/Q vssd1 vssd1 vccd1 vccd1 _09397_/C sky130_fd_sc_hd__or3_2
XFILLER_197_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_149_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_142_wb_clk_i clkbuf_5_26_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18317_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_145_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10170_ _10170_/A _10170_/B vssd1 vssd1 vccd1 vccd1 _10172_/C sky130_fd_sc_hd__xnor2_1
XFILLER_105_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_1363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_219_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13860_ _18829_/Q _13856_/X _13858_/X _18820_/Q _13859_/X vssd1 vssd1 vccd1 vccd1
+ _13860_/X sky130_fd_sc_hd__a221o_1
XFILLER_210_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12811_ _12533_/Y _17946_/Q _17951_/Q _12588_/B vssd1 vssd1 vccd1 vccd1 _12811_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_28_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13791_ _18288_/Q _13847_/A _13781_/X _18279_/Q vssd1 vssd1 vccd1 vccd1 _13791_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_43_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15530_ _15551_/A _16128_/B _15574_/C vssd1 vssd1 vccd1 vccd1 _15530_/X sky130_fd_sc_hd__or3_1
XTAP_1110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12742_ _12742_/A _12742_/B _12742_/C vssd1 vssd1 vccd1 vccd1 _12743_/C sky130_fd_sc_hd__and3_1
XFILLER_42_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15461_ _15460_/B _15458_/X _15460_/Y _15452_/X vssd1 vssd1 vccd1 vccd1 _18446_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_128_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12673_ _12672_/A _12672_/B _12537_/S vssd1 vssd1 vccd1 vccd1 _12673_/X sky130_fd_sc_hd__o21a_1
XFILLER_187_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_169_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_230_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17200_ _17213_/A _17200_/B vssd1 vssd1 vccd1 vccd1 _17200_/Y sky130_fd_sc_hd__nand2_1
X_11624_ _17857_/Q _11624_/B vssd1 vssd1 vccd1 vccd1 _11624_/X sky130_fd_sc_hd__or2_1
XTAP_1198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14412_ _17564_/A _14412_/B vssd1 vssd1 vccd1 vccd1 _14413_/A sky130_fd_sc_hd__and2_1
XFILLER_8_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18180_ _18184_/CLK _18180_/D vssd1 vssd1 vccd1 vccd1 _18180_/Q sky130_fd_sc_hd__dfxtp_1
X_15392_ _16909_/A vssd1 vssd1 vccd1 vccd1 _15993_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_204_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_168_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17131_ _17423_/A _17256_/C vssd1 vssd1 vccd1 vccd1 _17143_/B sky130_fd_sc_hd__nor2_2
XFILLER_50_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11555_ _17865_/Q vssd1 vssd1 vccd1 vccd1 _12261_/A sky130_fd_sc_hd__clkbuf_2
X_14343_ _18211_/Q _14305_/A _14342_/Y _14272_/A vssd1 vssd1 vccd1 vccd1 _14343_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_156_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10506_ _10443_/A _10503_/X _10505_/X vssd1 vssd1 vccd1 vccd1 _10506_/X sky130_fd_sc_hd__a21o_2
X_17062_ _17072_/A _17493_/B _17085_/C vssd1 vssd1 vccd1 vccd1 _17062_/X sky130_fd_sc_hd__or3_1
X_14274_ _14274_/A vssd1 vssd1 vccd1 vccd1 _18174_/D sky130_fd_sc_hd__clkbuf_1
X_11486_ _11719_/B _11364_/A _11257_/B _11595_/A vssd1 vssd1 vccd1 vccd1 _11486_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_7_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16013_ _16017_/B _16010_/X _16012_/Y _16008_/X vssd1 vssd1 vccd1 vccd1 _18580_/D
+ sky130_fd_sc_hd__o211a_1
X_13225_ _13233_/A _18068_/Q vssd1 vssd1 vccd1 vccd1 _13226_/A sky130_fd_sc_hd__and2_1
XFILLER_174_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10437_ _10456_/A _10441_/A vssd1 vssd1 vccd1 vccd1 _14289_/A sky130_fd_sc_hd__xor2_4
XFILLER_48_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_1274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13156_ _13164_/A _18037_/Q vssd1 vssd1 vccd1 vccd1 _13157_/A sky130_fd_sc_hd__and2_1
X_10368_ _09304_/A _09294_/B _09299_/C _09304_/C _10292_/S _10294_/X vssd1 vssd1 vccd1
+ vccd1 _10368_/X sky130_fd_sc_hd__mux4_1
XTAP_905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12107_ _12106_/A _12106_/B _13649_/A vssd1 vssd1 vccd1 vccd1 _12107_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_88_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_1288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13087_ _13094_/A vssd1 vssd1 vccd1 vccd1 _14377_/A sky130_fd_sc_hd__clkbuf_2
X_17964_ _17965_/CLK _17964_/D vssd1 vssd1 vccd1 vccd1 _17964_/Q sky130_fd_sc_hd__dfxtp_1
X_10299_ _09186_/B _09176_/B _09181_/C _09186_/C _09947_/A _10599_/S vssd1 vssd1 vccd1
+ vccd1 _10299_/X sky130_fd_sc_hd__mux4_1
X_16915_ _18830_/Q _18794_/Q _16925_/S vssd1 vssd1 vccd1 vccd1 _16915_/X sky130_fd_sc_hd__mux2_1
X_12038_ _12038_/A vssd1 vssd1 vccd1 vccd1 _13494_/B sky130_fd_sc_hd__buf_4
XFILLER_38_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17895_ _17895_/CLK _17895_/D vssd1 vssd1 vccd1 vccd1 _17895_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_66_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16846_ _18815_/Q _18779_/Q _16864_/S vssd1 vssd1 vccd1 vccd1 _16846_/X sky130_fd_sc_hd__mux2_1
XFILLER_65_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_207_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_225_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16777_ _16779_/B _16775_/X _16776_/Y _16760_/X vssd1 vssd1 vccd1 vccd1 _18763_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_53_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13989_ _18391_/Q _13666_/X _13986_/X _13988_/X vssd1 vssd1 vccd1 vccd1 _13989_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_34_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_206_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18516_ _18553_/CLK _18516_/D vssd1 vssd1 vccd1 vccd1 _18516_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_222_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15728_ _15730_/B _15726_/X _15727_/Y _15720_/X vssd1 vssd1 vccd1 vccd1 _18511_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_146_1302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_209_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_1204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_222_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18447_ _18473_/CLK _18447_/D vssd1 vssd1 vccd1 vccd1 _18447_/Q sky130_fd_sc_hd__dfxtp_1
X_15659_ _15661_/B _15657_/X _15658_/Y _15640_/X vssd1 vssd1 vccd1 vccd1 _18493_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_178_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09180_ _18605_/Q _18604_/Q _18603_/Q vssd1 vssd1 vccd1 vccd1 _09181_/D sky130_fd_sc_hd__or3_4
X_18378_ _18380_/CLK _18378_/D vssd1 vssd1 vccd1 vccd1 _18378_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_187_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17329_ _17471_/A _17399_/C vssd1 vssd1 vccd1 vccd1 _17336_/B sky130_fd_sc_hd__nor2_2
XFILLER_186_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_175_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_175_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_130_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08964_ _08966_/A vssd1 vssd1 vccd1 vccd1 _08964_/Y sky130_fd_sc_hd__inv_2
XFILLER_124_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_116_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_225_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09516_ _13416_/A _14386_/A _14383_/C _12217_/A vssd1 vssd1 vccd1 vccd1 _10990_/A
+ sky130_fd_sc_hd__o31a_4
XFILLER_225_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_227_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09447_ _09121_/A _09120_/Y _09222_/A _09446_/X vssd1 vssd1 vccd1 vccd1 _09447_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_73_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_223_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_227_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09378_ _18395_/Q _18394_/Q _18393_/Q vssd1 vssd1 vccd1 vccd1 _09381_/B sky130_fd_sc_hd__or3_4
XFILLER_40_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_185_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_166_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11340_ _11375_/A _11340_/B vssd1 vssd1 vccd1 vccd1 _11341_/A sky130_fd_sc_hd__and2_1
XFILLER_166_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11271_ _11315_/B _11268_/Y _11807_/A vssd1 vssd1 vccd1 vccd1 _11282_/B sky130_fd_sc_hd__a21oi_2
XFILLER_180_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19099__70 vssd1 vssd1 vccd1 vccd1 _19099__70/HI _19207_/A sky130_fd_sc_hd__conb_1
XFILLER_165_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13010_ _17992_/Q _12955_/A _13009_/Y _12721_/X _13007_/B vssd1 vssd1 vccd1 vccd1
+ _13010_/X sky130_fd_sc_hd__a221o_1
X_10222_ _10232_/A _10232_/B _10221_/X vssd1 vssd1 vccd1 vccd1 _10238_/B sky130_fd_sc_hd__a21o_1
XFILLER_180_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10153_ _10155_/A _10155_/C _10152_/X vssd1 vssd1 vccd1 vccd1 _10169_/A sky130_fd_sc_hd__o21ai_1
XTAP_5910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14961_ _14980_/A vssd1 vssd1 vccd1 vccd1 _14961_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_121_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10084_ _09287_/B _09282_/C _10096_/S vssd1 vssd1 vccd1 vccd1 _10084_/X sky130_fd_sc_hd__mux2_1
XTAP_5954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16700_ _16699_/B _16698_/X _16699_/Y _16683_/X vssd1 vssd1 vccd1 vccd1 _18743_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_102_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13912_ _18862_/Q _13596_/A _13561_/A _18865_/Q _13911_/X vssd1 vssd1 vccd1 vccd1
+ _13912_/X sky130_fd_sc_hd__a221o_1
XFILLER_43_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17680_ _17641_/X _17674_/Y _17675_/X _17676_/Y _18982_/Q vssd1 vssd1 vccd1 vccd1
+ _17681_/B sky130_fd_sc_hd__a32o_1
XTAP_5998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14892_ _15184_/A _14937_/B vssd1 vssd1 vccd1 vccd1 _14900_/B sky130_fd_sc_hd__nor2_1
XFILLER_207_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16631_ _16631_/A _16634_/B vssd1 vssd1 vccd1 vccd1 _16631_/Y sky130_fd_sc_hd__nand2_1
X_13843_ _18673_/Q _13842_/X _13546_/A _18670_/Q vssd1 vssd1 vccd1 vccd1 _13843_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_169_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16562_ _16575_/A _16562_/B vssd1 vssd1 vccd1 vccd1 _16562_/Y sky130_fd_sc_hd__nand2_1
X_13774_ _18648_/Q _13560_/A _13654_/X _18639_/Q _13773_/X vssd1 vssd1 vccd1 vccd1
+ _13774_/X sky130_fd_sc_hd__a221o_1
X_10986_ _14267_/A _09523_/X _10977_/X _10982_/X _10985_/X vssd1 vssd1 vccd1 vccd1
+ _19000_/D sky130_fd_sc_hd__a32o_1
X_18301_ _18307_/CLK _18301_/D vssd1 vssd1 vccd1 vccd1 _18301_/Q sky130_fd_sc_hd__dfxtp_1
X_15513_ _15962_/A _15548_/B vssd1 vssd1 vccd1 vccd1 _15525_/B sky130_fd_sc_hd__nor2_2
XFILLER_215_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_231_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_167_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12725_ _18089_/Q vssd1 vssd1 vccd1 vccd1 _12987_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_43_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16493_ _16493_/A vssd1 vssd1 vccd1 vccd1 _16509_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_71_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_206_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18232_ _18809_/CLK _18232_/D vssd1 vssd1 vccd1 vccd1 _18232_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_231_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15444_ _18479_/Q _18443_/Q _15458_/S vssd1 vssd1 vccd1 vccd1 _15444_/X sky130_fd_sc_hd__mux2_1
XFILLER_128_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12656_ _12656_/A _12656_/B vssd1 vssd1 vccd1 vccd1 _12656_/Y sky130_fd_sc_hd__nand2_1
XFILLER_141_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_230_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11607_ _12233_/A _17856_/Q _11624_/B vssd1 vssd1 vccd1 vccd1 _12235_/A sky130_fd_sc_hd__nand3_2
X_18163_ _18163_/CLK _18163_/D vssd1 vssd1 vccd1 vccd1 hold1/A sky130_fd_sc_hd__dfxtp_1
X_15375_ _15375_/A _15375_/B vssd1 vssd1 vccd1 vccd1 _15375_/Y sky130_fd_sc_hd__nand2_1
X_12587_ _12629_/A _17923_/Q vssd1 vssd1 vccd1 vccd1 _12590_/A sky130_fd_sc_hd__xnor2_1
XFILLER_15_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_209_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17114_ _18878_/Q _18842_/Q _17114_/S vssd1 vssd1 vccd1 vccd1 _17114_/X sky130_fd_sc_hd__mux2_1
XFILLER_172_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14326_ _14322_/Y _14325_/Y _14349_/A vssd1 vssd1 vccd1 vccd1 _14326_/X sky130_fd_sc_hd__mux2_1
X_18094_ _18094_/CLK _18094_/D vssd1 vssd1 vccd1 vccd1 _18094_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_7_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11538_ _11452_/A _11735_/B _11654_/C vssd1 vssd1 vccd1 vccd1 _11749_/A sky130_fd_sc_hd__a21oi_2
XFILLER_176_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17045_ _17168_/A vssd1 vssd1 vccd1 vccd1 _17091_/A sky130_fd_sc_hd__clkbuf_2
X_11469_ _11455_/D _11468_/X _11393_/X vssd1 vssd1 vccd1 vccd1 _11483_/B sky130_fd_sc_hd__o21ba_1
X_14257_ _14470_/B _14257_/B vssd1 vssd1 vccd1 vccd1 _14257_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_109_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13208_ _13208_/A _18061_/Q vssd1 vssd1 vccd1 vccd1 _13209_/A sky130_fd_sc_hd__and2_1
XFILLER_217_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14188_ _14188_/A vssd1 vssd1 vccd1 vccd1 _14330_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_174_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13139_ _13139_/A vssd1 vssd1 vccd1 vccd1 _18028_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_31_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18996_ _19000_/CLK _18996_/D vssd1 vssd1 vccd1 vccd1 _18996_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_112_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17947_ _17959_/CLK _17947_/D vssd1 vssd1 vccd1 vccd1 _17947_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_97_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_1277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_226_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17878_ _17884_/CLK _17878_/D vssd1 vssd1 vccd1 vccd1 _17878_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_65_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16829_ _16882_/A _16833_/B vssd1 vssd1 vccd1 vccd1 _16829_/Y sky130_fd_sc_hd__nand2_1
XFILLER_81_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_198_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09301_ _18500_/Q _18499_/Q _18498_/Q vssd1 vssd1 vccd1 vccd1 _09304_/B sky130_fd_sc_hd__or3_4
XFILLER_81_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_222_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_224_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09232_ _10826_/A _09232_/B _09232_/C _09232_/D vssd1 vssd1 vccd1 vccd1 _09238_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_179_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_222_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_222_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09163_ _18656_/Q _18655_/Q _18654_/Q vssd1 vssd1 vccd1 vccd1 _09165_/C sky130_fd_sc_hd__or3_4
XFILLER_119_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09094_ _18785_/Q _18784_/Q _18783_/Q vssd1 vssd1 vccd1 vccd1 _09098_/A sky130_fd_sc_hd__or3_4
XFILLER_119_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_135_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_1349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_89_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09996_ _09153_/B _10003_/S _09993_/X _10017_/S vssd1 vssd1 vccd1 vccd1 _09996_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_135_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08947_ _08948_/A vssd1 vssd1 vccd1 vccd1 _08947_/Y sky130_fd_sc_hd__inv_2
XTAP_4516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_218_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_229_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_218_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10840_ _09126_/A _09136_/B _09131_/A _09126_/D _10660_/X _10648_/X vssd1 vssd1 vccd1
+ vccd1 _10840_/X sky130_fd_sc_hd__mux4_2
XFILLER_72_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_226_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_198_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_213_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_1232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10771_ _09186_/A _09181_/A _09181_/D _09176_/D _10770_/X _10858_/S vssd1 vssd1 vccd1
+ vccd1 _10772_/C sky130_fd_sc_hd__mux4_2
XFILLER_53_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_201_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_213_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12510_ _12972_/A vssd1 vssd1 vccd1 vccd1 _12510_/X sky130_fd_sc_hd__buf_6
X_13490_ _13490_/A vssd1 vssd1 vccd1 vccd1 _13857_/A sky130_fd_sc_hd__buf_4
XFILLER_157_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_212_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12441_ _12441_/A vssd1 vssd1 vccd1 vccd1 _17901_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_12_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15160_ _15250_/A vssd1 vssd1 vccd1 vccd1 _15177_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_172_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12372_ _18989_/Q _18987_/Q vssd1 vssd1 vccd1 vccd1 _12381_/B sky130_fd_sc_hd__nor2_1
XFILLER_181_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14111_ _12042_/A _14103_/X _14110_/X _12027_/C vssd1 vssd1 vccd1 vccd1 _14111_/X
+ sky130_fd_sc_hd__a22o_1
X_11323_ _11323_/A _11323_/B _12299_/B vssd1 vssd1 vccd1 vccd1 _11323_/X sky130_fd_sc_hd__and3_1
X_15091_ _15115_/A _15094_/B vssd1 vssd1 vccd1 vccd1 _15091_/Y sky130_fd_sc_hd__nand2_1
XFILLER_5_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14042_ _18338_/Q _13575_/A _13576_/A _18329_/Q _14041_/X vssd1 vssd1 vccd1 vccd1
+ _14042_/X sky130_fd_sc_hd__a221o_2
X_11254_ _11653_/A _11730_/A vssd1 vssd1 vccd1 vccd1 _11254_/Y sky130_fd_sc_hd__nand2_1
XFILLER_109_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10205_ _10206_/A _10206_/B vssd1 vssd1 vccd1 vccd1 _10213_/B sky130_fd_sc_hd__xnor2_1
XFILLER_140_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18850_ _18866_/CLK _18850_/D vssd1 vssd1 vccd1 vccd1 _18850_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_192_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11185_ _17808_/Q _11185_/B vssd1 vssd1 vccd1 vccd1 _11186_/C sky130_fd_sc_hd__or2_1
X_17801_ _17851_/CLK _17801_/D vssd1 vssd1 vccd1 vccd1 _17801_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_121_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10136_ _19027_/Q _17980_/Q vssd1 vssd1 vccd1 vccd1 _10137_/B sky130_fd_sc_hd__or2_1
XFILLER_192_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18781_ _18821_/CLK _18781_/D vssd1 vssd1 vccd1 vccd1 _18781_/Q sky130_fd_sc_hd__dfxtp_4
XTAP_5740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15993_ _15993_/A _15993_/B vssd1 vssd1 vccd1 vccd1 _16003_/B sky130_fd_sc_hd__nor2_2
XTAP_5751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17732_ _17734_/A _19011_/Q vssd1 vssd1 vccd1 vccd1 _17733_/A sky130_fd_sc_hd__and2_1
XTAP_5773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14944_ _14944_/A vssd1 vssd1 vccd1 vccd1 _14992_/A sky130_fd_sc_hd__buf_2
X_10067_ _09657_/A _10045_/X _10053_/X _09720_/X _10066_/X vssd1 vssd1 vccd1 vccd1
+ _10068_/C sky130_fd_sc_hd__a32o_2
XFILLER_48_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17663_ _17663_/A _17663_/B vssd1 vssd1 vccd1 vccd1 _17663_/Y sky130_fd_sc_hd__nor2_1
X_14875_ _14875_/A _14875_/B vssd1 vssd1 vccd1 vccd1 _14875_/Y sky130_fd_sc_hd__nand2_1
XFILLER_21_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_223_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_224_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_103 _13858_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16614_ _18759_/Q _18723_/Q _16617_/S vssd1 vssd1 vccd1 vccd1 _16614_/X sky130_fd_sc_hd__mux2_1
XFILLER_165_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_223_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13826_ _18588_/Q _13759_/A _13780_/A _18579_/Q _13825_/X vssd1 vssd1 vccd1 vccd1
+ _13826_/X sky130_fd_sc_hd__a221o_1
XINSDIODE2_114 _15162_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17594_ _17610_/A _17594_/B vssd1 vssd1 vccd1 vccd1 _17595_/A sky130_fd_sc_hd__and2_1
XFILLER_189_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XINSDIODE2_125 _15257_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_1366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_223_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_136 _16566_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_91_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XINSDIODE2_147 input1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_1204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16545_ _16551_/B _16543_/X _16544_/X _16539_/X vssd1 vssd1 vccd1 vccd1 _18705_/D
+ sky130_fd_sc_hd__o211a_1
X_13757_ _18801_/Q _13617_/A _13730_/X _18804_/Q _13756_/X vssd1 vssd1 vccd1 vccd1
+ _13757_/X sky130_fd_sc_hd__a221o_2
XINSDIODE2_158 _18352_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_204_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10969_ _18227_/Q vssd1 vssd1 vccd1 vccd1 _14507_/A sky130_fd_sc_hd__clkbuf_2
XINSDIODE2_169 _18938_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_188_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_204_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12708_ _12708_/A _12708_/B _12707_/X vssd1 vssd1 vccd1 vccd1 _12709_/A sky130_fd_sc_hd__or3b_1
X_16476_ _16780_/A vssd1 vssd1 vccd1 vccd1 _16559_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_176_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13688_ _18606_/Q _13566_/A _13624_/A _18600_/Q _13687_/X vssd1 vssd1 vccd1 vccd1
+ _13688_/X sky130_fd_sc_hd__a221o_1
XFILLER_188_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18215_ _18217_/CLK _18215_/D vssd1 vssd1 vccd1 vccd1 _18215_/Q sky130_fd_sc_hd__dfxtp_1
X_15427_ _15739_/A vssd1 vssd1 vccd1 vccd1 _15516_/A sky130_fd_sc_hd__buf_2
X_19195_ _19195_/A _08996_/Y vssd1 vssd1 vccd1 vccd1 io_out[33] sky130_fd_sc_hd__ebufn_8
X_12639_ _12632_/A _12632_/B _12628_/A vssd1 vssd1 vccd1 vccd1 _12640_/B sky130_fd_sc_hd__o21ai_1
XFILLER_12_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18146_ _18147_/CLK _18146_/D vssd1 vssd1 vccd1 vccd1 _18146_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_15_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15358_ _15358_/A _15964_/B _15358_/C vssd1 vssd1 vccd1 vccd1 _15358_/X sky130_fd_sc_hd__or3_1
XFILLER_156_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14309_ _14319_/S _12131_/A _14307_/Y _14308_/X vssd1 vssd1 vccd1 vccd1 _14311_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_176_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18077_ _18085_/CLK _18077_/D vssd1 vssd1 vccd1 vccd1 _18077_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_89_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15289_ _17119_/A _17119_/B _16512_/C _15903_/C vssd1 vssd1 vccd1 vccd1 _15757_/A
+ sky130_fd_sc_hd__or4bb_4
XFILLER_172_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17028_ _17072_/A _17460_/B _17028_/C vssd1 vssd1 vccd1 vccd1 _17028_/X sky130_fd_sc_hd__or3_1
XFILLER_104_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09850_ _19028_/Q _12946_/A vssd1 vssd1 vccd1 vccd1 _09850_/X sky130_fd_sc_hd__and2_1
XFILLER_124_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09781_ _09781_/A _09781_/B vssd1 vssd1 vccd1 vccd1 _09781_/Y sky130_fd_sc_hd__nor2_1
XTAP_576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18979_ _18980_/CLK _18979_/D vssd1 vssd1 vccd1 vccd1 _18979_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_105_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_226_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_215_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_226_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_214_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_198_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_228_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_223_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_179_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_201_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_195_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_210_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09215_ _18671_/Q _18670_/Q _18669_/Q vssd1 vssd1 vccd1 vccd1 _09219_/A sky130_fd_sc_hd__or3_4
XFILLER_33_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09146_ _18704_/Q _18703_/Q _18702_/Q vssd1 vssd1 vccd1 vccd1 _09148_/C sky130_fd_sc_hd__or3_4
XFILLER_175_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09077_ _09083_/A _09081_/B _17831_/Q vssd1 vssd1 vccd1 vccd1 _09078_/A sky130_fd_sc_hd__and3_1
XFILLER_107_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_49_wb_clk_i clkbuf_5_16_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18823_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_155_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19069__40 vssd1 vssd1 vccd1 vccd1 _19069__40/HI _19163_/A sky130_fd_sc_hd__conb_1
XFILLER_162_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09979_ _09979_/A vssd1 vssd1 vccd1 vccd1 _12126_/A sky130_fd_sc_hd__buf_2
XTAP_5047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12990_ _12990_/A vssd1 vssd1 vccd1 vccd1 _12990_/Y sky130_fd_sc_hd__inv_2
XFILLER_183_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11941_ _11975_/A _11942_/A vssd1 vssd1 vccd1 vccd1 _13426_/A sky130_fd_sc_hd__xnor2_4
XFILLER_206_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_229_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_205_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_229_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14660_ _17663_/A _14660_/B vssd1 vssd1 vccd1 vccd1 _16932_/A sky130_fd_sc_hd__or2_4
XTAP_2933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11872_ _11879_/A _11872_/B vssd1 vssd1 vccd1 vccd1 _17829_/D sky130_fd_sc_hd__nor2_1
XFILLER_73_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13611_ _14014_/A vssd1 vssd1 vccd1 vccd1 _13612_/A sky130_fd_sc_hd__buf_6
XTAP_2977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10823_ _09237_/A _09227_/B _09232_/C _09237_/C _10695_/X _10852_/A vssd1 vssd1 vccd1
+ vccd1 _10823_/X sky130_fd_sc_hd__mux4_1
XFILLER_207_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14591_ _18174_/Q _18173_/Q _18170_/Q _18169_/Q vssd1 vssd1 vccd1 vccd1 _14609_/B
+ sky130_fd_sc_hd__or4bb_2
XTAP_2988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16330_ _16329_/B _16328_/X _16329_/Y _16314_/X vssd1 vssd1 vccd1 vccd1 _18653_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_186_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13542_ _13664_/A vssd1 vssd1 vccd1 vccd1 _13749_/A sky130_fd_sc_hd__buf_4
XFILLER_207_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10754_ _10763_/S vssd1 vssd1 vccd1 vccd1 _10877_/B sky130_fd_sc_hd__buf_4
XFILLER_200_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16261_ _16503_/A vssd1 vssd1 vccd1 vccd1 _16310_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_40_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13473_ _13480_/A _13473_/B vssd1 vssd1 vccd1 vccd1 _18159_/D sky130_fd_sc_hd__nor2_1
X_10685_ _10818_/B vssd1 vssd1 vccd1 vccd1 _10838_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_200_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18000_ _18088_/CLK _18000_/D vssd1 vssd1 vccd1 vccd1 _18000_/Q sky130_fd_sc_hd__dfxtp_1
X_15212_ _15220_/A _15371_/B _15257_/C vssd1 vssd1 vccd1 vccd1 _15212_/X sky130_fd_sc_hd__or3_1
XFILLER_12_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_185_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12424_ _12424_/A vssd1 vssd1 vccd1 vccd1 _17899_/D sky130_fd_sc_hd__clkbuf_1
X_16192_ _18657_/Q _18621_/Q _16192_/S vssd1 vssd1 vccd1 vccd1 _16192_/X sky130_fd_sc_hd__mux2_1
X_15143_ _15187_/A vssd1 vssd1 vccd1 vccd1 _15143_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_153_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12355_ _18991_/Q _12426_/C vssd1 vssd1 vccd1 vccd1 _12420_/B sky130_fd_sc_hd__nor2_1
XFILLER_86_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11306_ _11392_/B vssd1 vssd1 vccd1 vccd1 _11442_/A sky130_fd_sc_hd__clkbuf_2
X_15074_ _15218_/A _15085_/B vssd1 vssd1 vccd1 vccd1 _15082_/B sky130_fd_sc_hd__nor2_2
XFILLER_141_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12286_ _11530_/B _12272_/X _12284_/X _12285_/X vssd1 vssd1 vccd1 vccd1 _17871_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_99_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14025_ _18878_/Q _14015_/X _14018_/X _14024_/X vssd1 vssd1 vccd1 vccd1 _14025_/X
+ sky130_fd_sc_hd__a211o_2
X_11237_ _11892_/A _11237_/B _11237_/C vssd1 vssd1 vccd1 vccd1 _11242_/B sky130_fd_sc_hd__and3_1
X_18902_ _18902_/CLK _18902_/D vssd1 vssd1 vccd1 vccd1 _18902_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_206_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_214_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18833_ _18871_/CLK _18833_/D vssd1 vssd1 vccd1 vccd1 _18833_/Q sky130_fd_sc_hd__dfxtp_2
X_11168_ _17812_/Q _17811_/Q _17810_/Q _17809_/Q vssd1 vssd1 vccd1 vccd1 _11169_/C
+ sky130_fd_sc_hd__or4_1
XFILLER_150_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_228_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10119_ _10120_/A _10120_/B _10120_/C vssd1 vssd1 vccd1 vccd1 _10133_/A sky130_fd_sc_hd__a21oi_4
X_18764_ _18764_/CLK _18764_/D vssd1 vssd1 vccd1 vccd1 _18764_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_5570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15976_ _15984_/A _16128_/B _16021_/C vssd1 vssd1 vccd1 vccd1 _15976_/X sky130_fd_sc_hd__or3_1
X_11099_ _11099_/A vssd1 vssd1 vccd1 vccd1 _17794_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_83_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17715_ _17723_/A _19003_/Q vssd1 vssd1 vccd1 vccd1 _17716_/A sky130_fd_sc_hd__and2_1
XFILLER_76_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_222_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14927_ _18357_/Q _18321_/Q _14934_/S vssd1 vssd1 vccd1 vccd1 _14927_/X sky130_fd_sc_hd__mux2_1
XFILLER_110_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18695_ _18732_/CLK _18695_/D vssd1 vssd1 vccd1 vccd1 _18695_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_212_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17646_ _17645_/X _17635_/Y _17631_/X _17636_/Y _18974_/Q vssd1 vssd1 vccd1 vccd1
+ _17647_/B sky130_fd_sc_hd__a32o_1
XFILLER_110_1359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14858_ _14872_/A _14861_/B vssd1 vssd1 vccd1 vccd1 _14858_/Y sky130_fd_sc_hd__nand2_1
XFILLER_17_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_224_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13809_ _18405_/Q _13738_/A _13807_/X _13808_/X vssd1 vssd1 vccd1 vccd1 _13809_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_205_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17577_ _17576_/Y _17552_/A _14414_/A vssd1 vssd1 vccd1 vccd1 _17577_/Y sky130_fd_sc_hd__a21oi_1
X_14789_ _14788_/B _14787_/X _14788_/Y _14778_/X vssd1 vssd1 vccd1 vccd1 _18287_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_90_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_223_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_205_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16528_ _18138_/Q _16528_/B vssd1 vssd1 vccd1 vccd1 _16641_/A sky130_fd_sc_hd__nand2_2
XFILLER_189_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_220_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16459_ _16521_/A vssd1 vssd1 vccd1 vccd1 _16507_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_149_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09000_ _09003_/A vssd1 vssd1 vccd1 vccd1 _09000_/Y sky130_fd_sc_hd__inv_2
XFILLER_176_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19178_ _19178_/A _09010_/Y vssd1 vssd1 vccd1 vccd1 io_out[16] sky130_fd_sc_hd__ebufn_8
XFILLER_129_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18129_ _19028_/CLK _18129_/D vssd1 vssd1 vccd1 vccd1 _18129_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_118_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09902_ _09902_/A _09910_/B vssd1 vssd1 vccd1 vccd1 _10294_/A sky130_fd_sc_hd__or2b_2
XFILLER_104_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_1283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09833_ _09855_/A _09833_/B vssd1 vssd1 vccd1 vccd1 _12109_/B sky130_fd_sc_hd__xnor2_1
XFILLER_112_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09764_ _09764_/A _09764_/B vssd1 vssd1 vccd1 vccd1 _09792_/B sky130_fd_sc_hd__xnor2_1
XFILLER_230_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_167_wb_clk_i clkbuf_5_10_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18087_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_230_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09695_ _18248_/Q _18247_/Q _18246_/Q vssd1 vssd1 vccd1 vccd1 _09695_/X sky130_fd_sc_hd__or3_4
XFILLER_27_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_186_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_210_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_194_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10470_ _09237_/D _09232_/D _09227_/C _09232_/B _10464_/X _10235_/A vssd1 vssd1 vccd1
+ vccd1 _10470_/X sky130_fd_sc_hd__mux4_1
XFILLER_6_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09129_ _18812_/Q _18811_/Q _18810_/Q vssd1 vssd1 vccd1 vccd1 _09131_/C sky130_fd_sc_hd__or3_4
XFILLER_108_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12140_ _12158_/A _12169_/A vssd1 vssd1 vccd1 vccd1 _12141_/B sky130_fd_sc_hd__xor2_1
XFILLER_163_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12071_ _09692_/A _09719_/B _12070_/Y vssd1 vssd1 vccd1 vccd1 _12084_/A sky130_fd_sc_hd__a21oi_2
XFILLER_172_1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11022_ _13375_/C _11037_/C _13375_/B vssd1 vssd1 vccd1 vccd1 _11023_/A sky130_fd_sc_hd__and3b_1
XFILLER_110_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15830_ _18536_/Q _15829_/B _15829_/Y _15823_/X vssd1 vssd1 vccd1 vccd1 _18536_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_4110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15761_ _15892_/B vssd1 vssd1 vccd1 vccd1 _15811_/C sky130_fd_sc_hd__clkbuf_2
XTAP_4165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12973_ _12967_/A _12949_/Y _12971_/X _12972_/X vssd1 vssd1 vccd1 vccd1 _17975_/D
+ sky130_fd_sc_hd__a211o_1
XFILLER_45_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17500_ _18974_/Q _18938_/Q _17515_/S vssd1 vssd1 vccd1 vccd1 _17500_/X sky130_fd_sc_hd__mux2_1
XFILLER_206_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14712_ _18267_/Q _14715_/B _14711_/X _14692_/X vssd1 vssd1 vccd1 vccd1 _18267_/D
+ sky130_fd_sc_hd__o211a_1
X_18480_ _18482_/CLK _18480_/D vssd1 vssd1 vccd1 vccd1 _18480_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11924_ _11924_/A _12126_/B vssd1 vssd1 vccd1 vccd1 _11924_/Y sky130_fd_sc_hd__nand2_1
X_15692_ _15694_/B _15690_/X _15691_/Y _15681_/X vssd1 vssd1 vccd1 vccd1 _18502_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_3475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17431_ _18956_/Q _18920_/Q _17447_/S vssd1 vssd1 vccd1 vccd1 _17431_/X sky130_fd_sc_hd__mux2_1
XTAP_2752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14643_ _18252_/Q _14646_/B _14642_/X _14629_/X vssd1 vssd1 vccd1 vccd1 _18252_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_60_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11855_ _18156_/Q _11813_/Y _11853_/X _14185_/A vssd1 vssd1 vccd1 vccd1 _17827_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_72_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_198_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10806_ _10779_/X _10910_/D _10803_/X _10805_/X _10671_/B vssd1 vssd1 vccd1 vccd1
+ _10806_/X sky130_fd_sc_hd__a311o_1
XFILLER_60_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17362_ _17360_/B _17359_/X _17360_/Y _17361_/X vssd1 vssd1 vccd1 vccd1 _18902_/D
+ sky130_fd_sc_hd__o211a_1
X_14574_ _14606_/A _14574_/B vssd1 vssd1 vccd1 vccd1 _14574_/Y sky130_fd_sc_hd__nand2_1
XFILLER_92_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11786_ _11786_/A _11786_/B vssd1 vssd1 vccd1 vccd1 _11786_/Y sky130_fd_sc_hd__nand2_1
XFILLER_201_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16313_ _16325_/A _16317_/B vssd1 vssd1 vccd1 vccd1 _16313_/Y sky130_fd_sc_hd__nand2_1
XFILLER_198_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13525_ _13525_/A vssd1 vssd1 vccd1 vccd1 _13525_/X sky130_fd_sc_hd__buf_6
XFILLER_13_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10737_ _09098_/A _09103_/D _10737_/S vssd1 vssd1 vccd1 vccd1 _10738_/B sky130_fd_sc_hd__mux2_1
XFILLER_140_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17293_ _17331_/A vssd1 vssd1 vccd1 vccd1 _17351_/B sky130_fd_sc_hd__buf_2
XFILLER_201_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19032_ _19032_/CLK _19032_/D vssd1 vssd1 vccd1 vccd1 _19032_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16244_ _16243_/B _16242_/X _16243_/Y _16230_/X vssd1 vssd1 vccd1 vccd1 _18632_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_185_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13456_ _13458_/B _13456_/B _13456_/C vssd1 vssd1 vccd1 vccd1 _13457_/A sky130_fd_sc_hd__and3b_1
XFILLER_127_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10668_ _10668_/A vssd1 vssd1 vccd1 vccd1 _10811_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_12_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12407_ _12414_/B _12490_/A _12407_/C vssd1 vssd1 vccd1 vccd1 _12408_/A sky130_fd_sc_hd__and3b_1
X_16175_ _16202_/A _16175_/B vssd1 vssd1 vccd1 vccd1 _16175_/Y sky130_fd_sc_hd__nand2_1
XFILLER_177_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10599_ _09676_/X _09678_/X _10599_/S vssd1 vssd1 vccd1 vccd1 _10599_/X sky130_fd_sc_hd__mux2_1
XFILLER_127_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13387_ _18117_/Q _13386_/Y _13342_/X _13383_/A _11026_/X vssd1 vssd1 vccd1 vccd1
+ _18117_/D sky130_fd_sc_hd__o2111a_1
XFILLER_182_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_217_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15126_ _18406_/Q _18370_/Q _15141_/S vssd1 vssd1 vccd1 vccd1 _15126_/X sky130_fd_sc_hd__mux2_1
XFILLER_142_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12338_ _13153_/A _12338_/B vssd1 vssd1 vccd1 vccd1 _17885_/D sky130_fd_sc_hd__nor2_1
XFILLER_5_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15057_ _18388_/Q _18352_/Q _15081_/S vssd1 vssd1 vccd1 vccd1 _15057_/X sky130_fd_sc_hd__mux2_1
Xclkbuf_5_30_0_wb_clk_i clkbuf_5_31_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_5_30_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_2
X_12269_ _12269_/A _12269_/B _12269_/C vssd1 vssd1 vccd1 vccd1 _12269_/X sky130_fd_sc_hd__and3_1
XFILLER_218_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14008_ _12019_/A _13977_/X _13992_/X _14007_/X vssd1 vssd1 vccd1 vccd1 _14009_/D
+ sky130_fd_sc_hd__a211o_1
XFILLER_96_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18816_ _18826_/CLK _18816_/D vssd1 vssd1 vccd1 vccd1 _18816_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_83_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_228_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15959_ _16216_/A vssd1 vssd1 vccd1 vccd1 _16003_/A sky130_fd_sc_hd__clkbuf_2
X_18747_ _18752_/CLK _18747_/D vssd1 vssd1 vccd1 vccd1 _18747_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_95_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18678_ _18686_/CLK _18678_/D vssd1 vssd1 vccd1 vccd1 _18678_/Q sky130_fd_sc_hd__dfxtp_2
X_09480_ _09463_/X _09461_/A _09471_/B _18146_/D vssd1 vssd1 vccd1 vccd1 _18145_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_224_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_1333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17629_ _17638_/A _17629_/B vssd1 vssd1 vccd1 vccd1 _17630_/A sky130_fd_sc_hd__and2_1
XFILLER_211_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_225_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_180_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_195_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_1367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_219_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_219_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19039__10 vssd1 vssd1 vccd1 vccd1 _19039__10/HI _19133_/A sky130_fd_sc_hd__conb_1
XFILLER_28_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09816_ _09816_/A _09816_/B _09816_/C vssd1 vssd1 vccd1 vccd1 _09817_/A sky130_fd_sc_hd__and3_1
XFILLER_87_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_219_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09747_ _09748_/A _09753_/A _09748_/C vssd1 vssd1 vccd1 vccd1 _09749_/B sky130_fd_sc_hd__a21o_1
XFILLER_39_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_227_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09678_ _18245_/Q _18244_/Q _18243_/Q vssd1 vssd1 vccd1 vccd1 _09678_/X sky130_fd_sc_hd__or3_4
XTAP_2026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11640_ _17863_/Q _11668_/A vssd1 vssd1 vccd1 vccd1 _11640_/Y sky130_fd_sc_hd__nand2_1
XTAP_1369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_230_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_168_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11571_ _11549_/X _11565_/B _11570_/X _11563_/X vssd1 vssd1 vccd1 vccd1 _11571_/Y
+ sky130_fd_sc_hd__a31oi_1
XFILLER_196_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_64_wb_clk_i _18759_/CLK vssd1 vssd1 vccd1 vccd1 _18719_/CLK sky130_fd_sc_hd__clkbuf_16
X_13310_ _13310_/A _13310_/B _13310_/C vssd1 vssd1 vccd1 vccd1 _13311_/D sky130_fd_sc_hd__or3_1
XFILLER_195_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10522_ _10522_/A vssd1 vssd1 vccd1 vccd1 _10522_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_168_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14290_ _14187_/A _12065_/A _12100_/A _14237_/X _19000_/Q vssd1 vssd1 vccd1 vccd1
+ _14290_/X sky130_fd_sc_hd__a221o_1
XFILLER_161_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13241_ _13241_/A vssd1 vssd1 vccd1 vccd1 _18074_/D sky130_fd_sc_hd__clkbuf_1
X_10453_ _10443_/X _10447_/X _10452_/X _10270_/A vssd1 vssd1 vccd1 vccd1 _10453_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_170_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10384_ _09959_/X _10381_/X _10383_/X _10356_/A vssd1 vssd1 vccd1 vccd1 _10384_/X
+ sky130_fd_sc_hd__a211o_1
X_13172_ _13172_/A vssd1 vssd1 vccd1 vccd1 _18043_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_100_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12123_ _12123_/A _13526_/A vssd1 vssd1 vccd1 vccd1 _12123_/Y sky130_fd_sc_hd__nand2_1
X_17980_ _17990_/CLK _17980_/D vssd1 vssd1 vccd1 vccd1 _17980_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_97_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16931_ _16930_/B _16929_/X _16930_/Y _16917_/X vssd1 vssd1 vccd1 vccd1 _18797_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_117_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12054_ _12054_/A _12054_/B _12054_/C _12054_/D vssd1 vssd1 vccd1 vccd1 _12054_/X
+ sky130_fd_sc_hd__or4_1
XFILLER_133_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11005_ _17809_/Q vssd1 vssd1 vccd1 vccd1 _11190_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_120_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16862_ _16862_/A vssd1 vssd1 vccd1 vccd1 _17458_/A sky130_fd_sc_hd__buf_4
XFILLER_37_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18601_ _18635_/CLK _18601_/D vssd1 vssd1 vccd1 vccd1 _18601_/Q sky130_fd_sc_hd__dfxtp_4
X_15813_ _15863_/A vssd1 vssd1 vccd1 vccd1 _15838_/S sky130_fd_sc_hd__clkbuf_2
X_16793_ _16792_/B _16791_/X _16792_/Y _16781_/X vssd1 vssd1 vccd1 vccd1 _18767_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_203_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_219_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18532_ _18532_/CLK _18532_/D vssd1 vssd1 vccd1 vccd1 _18532_/Q sky130_fd_sc_hd__dfxtp_2
X_15744_ _15743_/B _15742_/X _15743_/Y _15740_/X vssd1 vssd1 vccd1 vccd1 _18515_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_3250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12956_ _12956_/A vssd1 vssd1 vccd1 vccd1 _12958_/B sky130_fd_sc_hd__inv_2
XTAP_3261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18463_ _18485_/CLK _18463_/D vssd1 vssd1 vccd1 vccd1 _18463_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11907_ _12141_/A vssd1 vssd1 vccd1 vccd1 _12171_/B sky130_fd_sc_hd__clkbuf_2
X_15675_ _16431_/A vssd1 vssd1 vccd1 vccd1 _16287_/A sky130_fd_sc_hd__buf_4
XTAP_2560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12887_ _17957_/Q _17958_/Q _12881_/B _17959_/Q vssd1 vssd1 vccd1 vccd1 _12888_/C
+ sky130_fd_sc_hd__a31o_1
XTAP_2571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17414_ _17536_/B vssd1 vssd1 vccd1 vccd1 _17460_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_14626_ _16886_/A vssd1 vssd1 vccd1 vccd1 _16889_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_60_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18394_ _18398_/CLK _18394_/D vssd1 vssd1 vccd1 vccd1 _18394_/Q sky130_fd_sc_hd__dfxtp_4
X_11838_ _11451_/Y _11835_/X _11837_/X _11491_/Y vssd1 vssd1 vccd1 vccd1 _11838_/X
+ sky130_fd_sc_hd__a211o_1
XTAP_1870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17345_ _17392_/A _17349_/B vssd1 vssd1 vccd1 vccd1 _17345_/Y sky130_fd_sc_hd__nand2_1
X_14557_ _14604_/A _14559_/B vssd1 vssd1 vccd1 vccd1 _14557_/Y sky130_fd_sc_hd__nand2_1
X_11769_ _11775_/A _11781_/B vssd1 vssd1 vccd1 vccd1 _11769_/X sky130_fd_sc_hd__or2_1
XFILLER_13_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_187_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13508_ _13508_/A vssd1 vssd1 vccd1 vccd1 _13508_/X sky130_fd_sc_hd__buf_6
XFILLER_144_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17276_ _18881_/Q _17275_/B _17275_/Y _17260_/X vssd1 vssd1 vccd1 vccd1 _18881_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_147_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14488_ _14488_/A vssd1 vssd1 vccd1 vccd1 _18218_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_228_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19015_ _19029_/CLK _19015_/D vssd1 vssd1 vccd1 vccd1 _19015_/Q sky130_fd_sc_hd__dfxtp_1
X_16227_ _16265_/A _16229_/B vssd1 vssd1 vccd1 vccd1 _16227_/Y sky130_fd_sc_hd__nand2_1
XFILLER_174_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13439_ _13439_/A _13439_/B vssd1 vssd1 vccd1 vccd1 _13439_/Y sky130_fd_sc_hd__nand2_1
XFILLER_220_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16158_ _16160_/B _16156_/X _16157_/Y _16139_/X vssd1 vssd1 vccd1 vccd1 _18613_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_161_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_154_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15109_ _15255_/A _15134_/B vssd1 vssd1 vccd1 vccd1 _15118_/B sky130_fd_sc_hd__nor2_1
XFILLER_114_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19123__94 vssd1 vssd1 vccd1 vccd1 _19123__94/HI _19231_/A sky130_fd_sc_hd__conb_1
X_08980_ _08998_/A vssd1 vssd1 vccd1 vccd1 _08985_/A sky130_fd_sc_hd__buf_12
X_16089_ _16115_/A _16692_/B _16115_/C vssd1 vssd1 vccd1 vccd1 _16089_/X sky130_fd_sc_hd__or3_1
XFILLER_142_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_228_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_217_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09601_ _09601_/A _09601_/B vssd1 vssd1 vccd1 vccd1 _09609_/A sky130_fd_sc_hd__or2_1
XFILLER_151_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09532_ _18108_/Q vssd1 vssd1 vccd1 vccd1 _09565_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_209_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_184_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09463_ _09463_/A vssd1 vssd1 vccd1 vccd1 _09463_/X sky130_fd_sc_hd__buf_2
XFILLER_52_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_225_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_224_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_225_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_145_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09394_ _18359_/Q _18358_/Q _18357_/Q vssd1 vssd1 vccd1 vccd1 _09397_/B sky130_fd_sc_hd__or3_2
XFILLER_52_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_212_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_149_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_195_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_191_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_182_wb_clk_i clkbuf_5_8_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _19026_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_154_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_111_wb_clk_i clkbuf_5_29_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18532_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_43_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_219_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12810_ _12806_/Y _12807_/X _12808_/X _12809_/Y vssd1 vssd1 vccd1 vccd1 _12813_/C
+ sky130_fd_sc_hd__a22o_1
X_13790_ _12042_/A _13779_/X _13789_/X _12028_/D vssd1 vssd1 vccd1 vccd1 _13829_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_16_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12741_ _19012_/Q _19011_/Q _19014_/Q _19013_/Q vssd1 vssd1 vccd1 vccd1 _12742_/C
+ sky130_fd_sc_hd__and4_1
XFILLER_203_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15460_ _15511_/A _15460_/B vssd1 vssd1 vccd1 vccd1 _15460_/Y sky130_fd_sc_hd__nand2_1
XTAP_1155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_230_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12672_ _12672_/A _12672_/B vssd1 vssd1 vccd1 vccd1 _12672_/Y sky130_fd_sc_hd__nand2_1
XTAP_1166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14411_ _14414_/B _14386_/Y _14410_/X _18193_/Q vssd1 vssd1 vccd1 vccd1 _14412_/B
+ sky130_fd_sc_hd__a22o_1
X_11623_ _11689_/A _11623_/B vssd1 vssd1 vccd1 vccd1 _11623_/Y sky130_fd_sc_hd__nand2_1
XTAP_1199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15391_ _15390_/B _15388_/X _15390_/Y _15382_/X vssd1 vssd1 vccd1 vccd1 _18431_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_168_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17130_ _18845_/Q _17129_/B _17129_/Y _17117_/X vssd1 vssd1 vccd1 vccd1 _18845_/D
+ sky130_fd_sc_hd__o211a_1
X_14342_ _14342_/A _14342_/B vssd1 vssd1 vccd1 vccd1 _14342_/Y sky130_fd_sc_hd__nand2_1
X_11554_ _12267_/A _11339_/B _11553_/Y vssd1 vssd1 vccd1 vccd1 _11554_/X sky130_fd_sc_hd__a21o_1
XFILLER_195_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10505_ _10183_/A _10504_/X _10430_/X vssd1 vssd1 vccd1 vccd1 _10505_/X sky130_fd_sc_hd__a21bo_1
X_17061_ _18864_/Q _18828_/Q _17074_/S vssd1 vssd1 vccd1 vccd1 _17061_/X sky130_fd_sc_hd__mux2_1
XFILLER_6_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14273_ _14272_/X _14457_/B _18174_/Q _14463_/A vssd1 vssd1 vccd1 vccd1 _14274_/A
+ sky130_fd_sc_hd__and4b_1
X_11485_ _11455_/X _11465_/Y _11470_/Y _11476_/Y _11484_/X vssd1 vssd1 vccd1 vccd1
+ _11485_/X sky130_fd_sc_hd__a221o_1
XFILLER_10_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16012_ _16062_/A _16017_/B vssd1 vssd1 vccd1 vccd1 _16012_/Y sky130_fd_sc_hd__nand2_1
X_13224_ _13257_/A vssd1 vssd1 vccd1 vccd1 _13233_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_139_1310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10436_ _14307_/A _10939_/C _10436_/C vssd1 vssd1 vccd1 vccd1 _10436_/Y sky130_fd_sc_hd__nand3_1
XFILLER_48_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13155_ _13199_/A vssd1 vssd1 vccd1 vccd1 _13164_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_87_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10367_ _09294_/C _09299_/B _09304_/D _09299_/D _09950_/X _09959_/X vssd1 vssd1 vccd1
+ vccd1 _10367_/X sky130_fd_sc_hd__mux4_1
XTAP_906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12106_ _12106_/A _12106_/B _13649_/A vssd1 vssd1 vccd1 vccd1 _12106_/X sky130_fd_sc_hd__or3_1
XFILLER_3_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_215_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10298_ _10600_/A vssd1 vssd1 vccd1 vccd1 _10599_/S sky130_fd_sc_hd__buf_4
XTAP_939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13086_ _13086_/A vssd1 vssd1 vccd1 vccd1 _18005_/D sky130_fd_sc_hd__clkbuf_1
X_17963_ _17965_/CLK _17963_/D vssd1 vssd1 vccd1 vccd1 _17963_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_97_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_214_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16914_ _16916_/B _16912_/X _16913_/Y _16893_/X vssd1 vssd1 vccd1 vccd1 _18793_/D
+ sky130_fd_sc_hd__o211a_1
X_12037_ _12037_/A _12037_/B vssd1 vssd1 vccd1 vccd1 _12038_/A sky130_fd_sc_hd__and2_2
XFILLER_211_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17894_ _18989_/CLK _17894_/D vssd1 vssd1 vccd1 vccd1 _17894_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_226_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16845_ _16928_/A vssd1 vssd1 vccd1 vccd1 _16864_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_66_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16776_ _16813_/A _16779_/B vssd1 vssd1 vccd1 vccd1 _16776_/Y sky130_fd_sc_hd__nand2_1
XFILLER_230_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_225_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13988_ _18379_/Q _13719_/A _13721_/A _18403_/Q _13987_/X vssd1 vssd1 vccd1 vccd1
+ _13988_/X sky130_fd_sc_hd__a221o_1
XFILLER_18_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15727_ _15751_/A _15730_/B vssd1 vssd1 vccd1 vccd1 _15727_/Y sky130_fd_sc_hd__nand2_1
X_18515_ _18553_/CLK _18515_/D vssd1 vssd1 vccd1 vccd1 _18515_/Q sky130_fd_sc_hd__dfxtp_1
X_12939_ _12939_/A _12939_/B vssd1 vssd1 vccd1 vccd1 _17971_/D sky130_fd_sc_hd__nor2_1
XTAP_3080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15658_ _15691_/A _15661_/B vssd1 vssd1 vccd1 vccd1 _15658_/Y sky130_fd_sc_hd__nand2_1
X_18446_ _18448_/CLK _18446_/D vssd1 vssd1 vccd1 vccd1 _18446_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_222_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_146_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14609_ _14685_/B _14609_/B vssd1 vssd1 vccd1 vccd1 _14915_/A sky130_fd_sc_hd__or2_4
X_18377_ _18408_/CLK _18377_/D vssd1 vssd1 vccd1 vccd1 _18377_/Q sky130_fd_sc_hd__dfxtp_1
X_15589_ _15589_/A vssd1 vssd1 vccd1 vccd1 _15604_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_147_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17328_ _17327_/B _17326_/X _17327_/Y _17324_/X vssd1 vssd1 vccd1 vccd1 _18893_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_147_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17259_ _17273_/A _17263_/B vssd1 vssd1 vccd1 vccd1 _17259_/Y sky130_fd_sc_hd__nand2_1
XFILLER_135_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_216_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08963_ _08966_/A vssd1 vssd1 vccd1 vccd1 _08963_/Y sky130_fd_sc_hd__inv_2
XFILLER_69_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_229_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_190_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_217_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_112_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_225_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09515_ _17940_/Q _14510_/B vssd1 vssd1 vccd1 vccd1 _14383_/C sky130_fd_sc_hd__or2_4
XFILLER_37_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_197_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09446_ _09222_/B _09444_/Y _09445_/Y vssd1 vssd1 vccd1 vccd1 _09446_/X sky130_fd_sc_hd__a21o_1
XFILLER_25_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_227_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09377_ _18410_/Q _18409_/Q _18408_/Q vssd1 vssd1 vccd1 vccd1 _09381_/A sky130_fd_sc_hd__or3_4
XFILLER_12_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_197_1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_138_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11270_ _11368_/A _11926_/B _11334_/A vssd1 vssd1 vccd1 vccd1 _11807_/A sky130_fd_sc_hd__or3b_1
XFILLER_197_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10221_ _10220_/B _10221_/B vssd1 vssd1 vccd1 vccd1 _10221_/X sky130_fd_sc_hd__and2b_1
XFILLER_106_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10152_ _10155_/A _10155_/C _13389_/A vssd1 vssd1 vccd1 vccd1 _10152_/X sky130_fd_sc_hd__a21o_1
XFILLER_79_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14960_ _14995_/A _14960_/B vssd1 vssd1 vccd1 vccd1 _14960_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10083_ _09282_/A _09287_/C _10096_/S vssd1 vssd1 vccd1 vccd1 _10083_/X sky130_fd_sc_hd__mux2_1
XTAP_5944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_181_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13911_ _18859_/Q _13566_/A _13909_/X _13910_/X vssd1 vssd1 vccd1 vccd1 _13911_/X
+ sky130_fd_sc_hd__a211o_1
XTAP_5977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14891_ _14890_/B _14888_/X _14890_/Y _14881_/X vssd1 vssd1 vccd1 vccd1 _18311_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_47_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16630_ _18763_/Q _18727_/Q _16637_/S vssd1 vssd1 vccd1 vccd1 _16630_/X sky130_fd_sc_hd__mux2_1
X_13842_ _13842_/A vssd1 vssd1 vccd1 vccd1 _13842_/X sky130_fd_sc_hd__buf_6
XFILLER_210_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16561_ _18746_/Q _18710_/Q _16565_/S vssd1 vssd1 vccd1 vccd1 _16561_/X sky130_fd_sc_hd__mux2_1
X_13773_ _18642_/Q _13772_/X _13752_/X _18636_/Q vssd1 vssd1 vccd1 vccd1 _13773_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_15_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10985_ _14317_/A vssd1 vssd1 vccd1 vccd1 _10985_/X sky130_fd_sc_hd__clkbuf_2
X_15512_ _15511_/B _15510_/X _15511_/Y _15496_/X vssd1 vssd1 vccd1 vccd1 _18458_/D
+ sky130_fd_sc_hd__o211a_1
X_18300_ _18307_/CLK _18300_/D vssd1 vssd1 vccd1 vccd1 _18300_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_71_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12724_ _18153_/Q _12925_/B _12781_/B _18152_/Q vssd1 vssd1 vccd1 vccd1 _13271_/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_215_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16492_ _16499_/B _16490_/X _16491_/X _16477_/X vssd1 vssd1 vccd1 vccd1 _18693_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_167_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_230_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_230_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18231_ _18809_/CLK _18231_/D vssd1 vssd1 vccd1 vccd1 _18231_/Q sky130_fd_sc_hd__dfxtp_1
X_15443_ _15445_/B _15441_/X _15442_/Y _15428_/X vssd1 vssd1 vccd1 vccd1 _18442_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_54_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12655_ _12649_/A _12649_/B _12647_/A vssd1 vssd1 vccd1 vccd1 _12656_/B sky130_fd_sc_hd__a21o_1
XFILLER_231_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11606_ _17856_/Q _11624_/B vssd1 vssd1 vccd1 vccd1 _11606_/X sky130_fd_sc_hd__or2_1
X_18162_ _18163_/CLK _18162_/D vssd1 vssd1 vccd1 vccd1 _18162_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_90_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15374_ _18427_/Q _15375_/B _15373_/Y _15363_/X vssd1 vssd1 vccd1 vccd1 _18427_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_141_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12586_ _17926_/Q vssd1 vssd1 vccd1 vccd1 _12629_/A sky130_fd_sc_hd__buf_2
X_17113_ _17115_/B _17111_/X _17112_/Y _17096_/X vssd1 vssd1 vccd1 vccd1 _18841_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_11_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14325_ _14325_/A _14325_/B vssd1 vssd1 vccd1 vccd1 _14325_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_89_1326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18093_ _18095_/CLK _18093_/D vssd1 vssd1 vccd1 vccd1 _18093_/Q sky130_fd_sc_hd__dfxtp_1
X_11537_ _11513_/Y _11536_/X _11501_/X vssd1 vssd1 vccd1 vccd1 _11537_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_8_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17044_ _18823_/Q _17046_/B _17043_/Y _17040_/X vssd1 vssd1 vccd1 vccd1 _18823_/D
+ sky130_fd_sc_hd__o211a_1
X_14256_ _18209_/Q vssd1 vssd1 vccd1 vccd1 _14470_/B sky130_fd_sc_hd__clkbuf_2
X_11468_ _11365_/B _11468_/B _11539_/B vssd1 vssd1 vccd1 vccd1 _11468_/X sky130_fd_sc_hd__and3b_1
XFILLER_7_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13207_ _13207_/A vssd1 vssd1 vccd1 vccd1 _18059_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_124_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10419_ _10419_/A _10419_/B vssd1 vssd1 vccd1 vccd1 _10419_/Y sky130_fd_sc_hd__nand2_1
XFILLER_140_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14187_ _14187_/A _14204_/B vssd1 vssd1 vccd1 vccd1 _14188_/A sky130_fd_sc_hd__or2_1
X_11399_ _11399_/A vssd1 vssd1 vccd1 vccd1 _11413_/A sky130_fd_sc_hd__inv_2
XFILLER_112_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_225_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_217_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13138_ _13140_/A _18029_/Q vssd1 vssd1 vccd1 vccd1 _13139_/A sky130_fd_sc_hd__and2_1
XTAP_725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18995_ _19000_/CLK _18995_/D vssd1 vssd1 vccd1 vccd1 _18995_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13069_ _18000_/Q _12951_/A _13069_/S vssd1 vssd1 vccd1 vccd1 _13070_/B sky130_fd_sc_hd__mux2_1
X_17946_ _17965_/CLK _17946_/D vssd1 vssd1 vccd1 vccd1 _17946_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_24_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17877_ _17888_/CLK _17877_/D vssd1 vssd1 vccd1 vccd1 _17877_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16828_ _16828_/A vssd1 vssd1 vccd1 vccd1 _16882_/A sky130_fd_sc_hd__buf_2
XFILLER_81_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16759_ _16796_/A _16759_/B _16773_/C vssd1 vssd1 vccd1 vccd1 _16759_/X sky130_fd_sc_hd__or3_1
XFILLER_207_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09300_ _18497_/Q _18496_/Q _18495_/Q vssd1 vssd1 vccd1 vccd1 _09304_/A sky130_fd_sc_hd__or3_2
XFILLER_59_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_185_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_222_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09231_ _18941_/Q _18940_/Q _18939_/Q vssd1 vssd1 vccd1 vccd1 _09232_/D sky130_fd_sc_hd__or3_2
X_18429_ _18432_/CLK _18429_/D vssd1 vssd1 vccd1 vccd1 _18429_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_22_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_222_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09162_ _18629_/Q _18628_/Q _18627_/Q vssd1 vssd1 vccd1 vccd1 _10308_/A sky130_fd_sc_hd__or3_4
XFILLER_159_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_222_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_120_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09093_ _09093_/A _09093_/B _09093_/C _09093_/D vssd1 vssd1 vccd1 vccd1 _09104_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_135_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09995_ _09995_/A vssd1 vssd1 vccd1 vccd1 _10017_/S sky130_fd_sc_hd__buf_4
XTAP_5207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08946_ _08948_/A vssd1 vssd1 vccd1 vccd1 _08946_/Y sky130_fd_sc_hd__inv_2
XFILLER_130_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_218_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_218_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_226_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_213_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10770_ _10770_/A vssd1 vssd1 vccd1 vccd1 _10770_/X sky130_fd_sc_hd__buf_4
XFILLER_197_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_212_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09429_ _09429_/A vssd1 vssd1 vccd1 vccd1 _09430_/C sky130_fd_sc_hd__inv_2
XFILLER_40_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_200_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_1288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12440_ _12438_/Y _12440_/B _12467_/C vssd1 vssd1 vccd1 vccd1 _12441_/A sky130_fd_sc_hd__and3b_1
XFILLER_12_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_226_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12371_ _12467_/C vssd1 vssd1 vccd1 vccd1 _12459_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_154_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14110_ _18803_/Q _13838_/X _13575_/X _18806_/Q _14109_/X vssd1 vssd1 vccd1 vccd1
+ _14110_/X sky130_fd_sc_hd__a221o_2
XFILLER_153_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11322_ _17875_/Q vssd1 vssd1 vccd1 vccd1 _12299_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_176_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15090_ _18397_/Q _18361_/Q _15100_/S vssd1 vssd1 vccd1 vccd1 _15090_/X sky130_fd_sc_hd__mux2_1
XFILLER_180_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14041_ _18311_/Q _13619_/A _14037_/X _14040_/X vssd1 vssd1 vccd1 vccd1 _14041_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_10_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11253_ _11253_/A _11396_/B vssd1 vssd1 vccd1 vccd1 _11730_/A sky130_fd_sc_hd__nand2_1
XFILLER_84_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_1340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10204_ _10204_/A _10204_/B vssd1 vssd1 vccd1 vccd1 _10206_/B sky130_fd_sc_hd__xnor2_2
XFILLER_121_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11184_ _17808_/Q _17807_/Q _11184_/C vssd1 vssd1 vccd1 vccd1 _11196_/D sky130_fd_sc_hd__and3_1
XFILLER_121_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_192_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17800_ _17851_/CLK _17800_/D vssd1 vssd1 vccd1 vccd1 _17800_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_121_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10135_ _19027_/Q _17980_/Q vssd1 vssd1 vccd1 vccd1 _10135_/X sky130_fd_sc_hd__and2_1
X_15992_ _15991_/B _15990_/X _15991_/Y _15988_/X vssd1 vssd1 vccd1 vccd1 _18575_/D
+ sky130_fd_sc_hd__o211a_1
X_18780_ _18785_/CLK _18780_/D vssd1 vssd1 vccd1 vccd1 _18780_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_5730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14943_ _18361_/Q _18325_/Q _14955_/S vssd1 vssd1 vccd1 vccd1 _14943_/X sky130_fd_sc_hd__mux2_1
X_10066_ _10942_/A _10058_/X _10059_/X _10895_/A _10065_/X vssd1 vssd1 vccd1 vccd1
+ _10066_/X sky130_fd_sc_hd__a221o_1
X_17731_ _17731_/A vssd1 vssd1 vccd1 vccd1 _19009_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_94_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14874_ _18344_/Q _18308_/Q _14883_/S vssd1 vssd1 vccd1 vccd1 _14874_/X sky130_fd_sc_hd__mux2_1
XFILLER_1_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17662_ _17736_/A vssd1 vssd1 vccd1 vccd1 _17681_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_208_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_224_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_1262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_217_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16613_ _16757_/A _16650_/B vssd1 vssd1 vccd1 vccd1 _16623_/B sky130_fd_sc_hd__nor2_1
X_13825_ _18561_/Q _13664_/X _13821_/X _13824_/X vssd1 vssd1 vccd1 vccd1 _13825_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_217_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XINSDIODE2_104 _13858_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_169_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17593_ _17575_/X _17590_/Y _17582_/X _17592_/Y _18960_/Q vssd1 vssd1 vccd1 vccd1
+ _17594_/B sky130_fd_sc_hd__a32o_1
XFILLER_91_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_115 _15162_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_223_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XINSDIODE2_126 _15268_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_137 _15909_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16544_ _16555_/A _16692_/B _16568_/C vssd1 vssd1 vccd1 vccd1 _16544_/X sky130_fd_sc_hd__or3_1
XFILLER_90_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_148 input1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13756_ _18777_/Q _13749_/X _13751_/X _13755_/X vssd1 vssd1 vccd1 vccd1 _13756_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_204_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINSDIODE2_159 _18352_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_1216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10968_ _13411_/A _13411_/B _13411_/C _13411_/D vssd1 vssd1 vccd1 vccd1 _13415_/B
+ sky130_fd_sc_hd__or4_2
XFILLER_206_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_231_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12707_ _12707_/A _12707_/B _12707_/C vssd1 vssd1 vccd1 vccd1 _12707_/X sky130_fd_sc_hd__or3_1
X_16475_ _16510_/A _16475_/B vssd1 vssd1 vccd1 vccd1 _16475_/Y sky130_fd_sc_hd__nand2_1
XFILLER_43_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13687_ _18612_/Q _13559_/A _13490_/A _18603_/Q vssd1 vssd1 vccd1 vccd1 _13687_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_206_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10899_ _10899_/A _10899_/B vssd1 vssd1 vccd1 vccd1 _10899_/X sky130_fd_sc_hd__and2_1
XFILLER_176_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15426_ _15442_/A _15431_/B vssd1 vssd1 vccd1 vccd1 _15426_/Y sky130_fd_sc_hd__nand2_1
XFILLER_19_1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18214_ _18217_/CLK _18214_/D vssd1 vssd1 vccd1 vccd1 _18214_/Q sky130_fd_sc_hd__dfxtp_1
X_19194_ _19194_/A _08995_/Y vssd1 vssd1 vccd1 vccd1 io_out[32] sky130_fd_sc_hd__ebufn_8
X_12638_ _12638_/A _12638_/B vssd1 vssd1 vccd1 vccd1 _12640_/A sky130_fd_sc_hd__nor2_1
XFILLER_157_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_180_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15357_ _16865_/A vssd1 vssd1 vccd1 vccd1 _15964_/B sky130_fd_sc_hd__clkbuf_4
X_18145_ _18147_/CLK _18145_/D vssd1 vssd1 vccd1 vccd1 _18145_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_156_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_214_wb_clk_i clkbuf_5_9_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17817_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_200_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12569_ _12569_/A vssd1 vssd1 vccd1 vccd1 _12569_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_200_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14308_ _14187_/A _12063_/A _12102_/A _14237_/X _19000_/Q vssd1 vssd1 vccd1 vccd1
+ _14308_/X sky130_fd_sc_hd__a221o_1
X_18076_ _18085_/CLK _18076_/D vssd1 vssd1 vccd1 vccd1 _18076_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_172_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15288_ _15607_/C _15463_/B _15607_/B vssd1 vssd1 vccd1 vccd1 _17120_/A sky130_fd_sc_hd__nand3_4
XFILLER_85_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17027_ _17148_/A vssd1 vssd1 vccd1 vccd1 _17072_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_172_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14239_ _10236_/X _14205_/X _14238_/X vssd1 vssd1 vccd1 vccd1 _14239_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_171_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_217_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09780_ _10213_/A _09780_/B vssd1 vssd1 vccd1 vccd1 _09780_/Y sky130_fd_sc_hd__nand2_1
XFILLER_100_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18978_ _18980_/CLK _18978_/D vssd1 vssd1 vccd1 vccd1 _18978_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_85_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17929_ _17929_/CLK _17929_/D vssd1 vssd1 vccd1 vccd1 _17929_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_226_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_227_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_215_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_226_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_228_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_224_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_228_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_223_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_222_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_224_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09214_ _09214_/A _09214_/B _09214_/C _09214_/D vssd1 vssd1 vccd1 vccd1 _09220_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_195_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09145_ _18719_/Q _18718_/Q _18717_/Q vssd1 vssd1 vccd1 vccd1 _09148_/B sky130_fd_sc_hd__or3_4
XFILLER_136_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_136_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_159_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09076_ _09076_/A vssd1 vssd1 vccd1 vccd1 _19184_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_194_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_200_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09978_ _09921_/X _09941_/X _09956_/X _09966_/X _09977_/X vssd1 vssd1 vccd1 vccd1
+ _09978_/X sky130_fd_sc_hd__a2111o_1
XTAP_5037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19084__55 vssd1 vssd1 vccd1 vccd1 _19084__55/HI _19192_/A sky130_fd_sc_hd__conb_1
XFILLER_76_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_218_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_18_wb_clk_i clkbuf_5_5_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18870_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_5059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08929_ _09053_/A vssd1 vssd1 vccd1 vccd1 _11018_/A sky130_fd_sc_hd__buf_12
XTAP_4325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11940_ _11983_/A _11983_/B vssd1 vssd1 vccd1 vccd1 _12025_/B sky130_fd_sc_hd__nand2_1
XFILLER_85_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11871_ _18162_/Q _11867_/X _11870_/Y vssd1 vssd1 vccd1 vccd1 _11872_/B sky130_fd_sc_hd__a21oi_1
XTAP_2934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13610_ _12027_/B _13602_/X _13609_/X _13434_/C vssd1 vssd1 vccd1 vccd1 _13610_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_72_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10822_ _10822_/A _10822_/B _10822_/C _14330_/A vssd1 vssd1 vccd1 vccd1 _10822_/X
+ sky130_fd_sc_hd__or4b_1
X_14590_ _18242_/Q _14589_/B _14589_/Y _14587_/X vssd1 vssd1 vccd1 vccd1 _18242_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_32_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_164_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_207_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13541_ _13547_/B _13541_/B vssd1 vssd1 vccd1 vccd1 _13664_/A sky130_fd_sc_hd__nor2_1
XFILLER_25_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10753_ _10753_/A vssd1 vssd1 vccd1 vccd1 _10757_/A sky130_fd_sc_hd__buf_2
XFILLER_213_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16260_ _16566_/A vssd1 vssd1 vccd1 vccd1 _16503_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_125_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_185_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13472_ _17844_/Q _13457_/X _13465_/X vssd1 vssd1 vccd1 vccd1 _13473_/B sky130_fd_sc_hd__a21oi_1
XFILLER_41_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10684_ _09282_/A _09287_/B _09287_/C _09282_/C _10824_/A _10680_/A vssd1 vssd1 vccd1
+ vccd1 _10684_/X sky130_fd_sc_hd__mux4_1
XFILLER_201_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15211_ _15211_/A vssd1 vssd1 vccd1 vccd1 _15257_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_16_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12423_ _12459_/A _12423_/B _12430_/B vssd1 vssd1 vccd1 vccd1 _12424_/A sky130_fd_sc_hd__and3_1
XFILLER_200_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16191_ _16783_/A _16205_/B vssd1 vssd1 vccd1 vccd1 _16202_/B sky130_fd_sc_hd__nor2_2
XFILLER_166_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15142_ _15182_/A _15142_/B vssd1 vssd1 vccd1 vccd1 _15142_/Y sky130_fd_sc_hd__nand2_1
X_12354_ _18106_/Q _18990_/Q _12401_/B vssd1 vssd1 vccd1 vccd1 _12426_/C sky130_fd_sc_hd__or3_1
XFILLER_5_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11305_ _13501_/A _11392_/B vssd1 vssd1 vccd1 vccd1 _11305_/X sky130_fd_sc_hd__or2_1
X_15073_ _18356_/Q _15072_/B _15072_/Y _15066_/X vssd1 vssd1 vccd1 vccd1 _18356_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_99_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12285_ _12285_/A _12285_/B _12285_/C vssd1 vssd1 vccd1 vccd1 _12285_/X sky130_fd_sc_hd__and3_1
XFILLER_4_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_5_20_0_wb_clk_i clkbuf_5_21_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_5_20_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_2
X_14024_ _18863_/Q _13525_/X _13621_/X _18866_/Q _14023_/X vssd1 vssd1 vccd1 vccd1
+ _14024_/X sky130_fd_sc_hd__a221o_1
X_18901_ _18902_/CLK _18901_/D vssd1 vssd1 vccd1 vccd1 _18901_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_141_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11236_ _11001_/C _11234_/A _11235_/Y vssd1 vssd1 vccd1 vccd1 _17821_/D sky130_fd_sc_hd__a21oi_1
XFILLER_49_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_106_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_214_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18832_ _18849_/CLK _18832_/D vssd1 vssd1 vccd1 vccd1 _18832_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_95_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11167_ _11181_/A _17805_/Q vssd1 vssd1 vccd1 vccd1 _11169_/B sky130_fd_sc_hd__nand2_1
XFILLER_67_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10118_ _18127_/Q _10118_/B vssd1 vssd1 vccd1 vccd1 _10120_/C sky130_fd_sc_hd__xnor2_1
X_18763_ _18799_/CLK _18763_/D vssd1 vssd1 vccd1 vccd1 _18763_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_121_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15975_ _15975_/A vssd1 vssd1 vccd1 vccd1 _16021_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_48_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11098_ _11281_/A _17824_/Q _11113_/S vssd1 vssd1 vccd1 vccd1 _11099_/A sky130_fd_sc_hd__mux2_1
XFILLER_95_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17714_ _17736_/A vssd1 vssd1 vccd1 vccd1 _17723_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_208_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14926_ _15218_/A _14937_/B vssd1 vssd1 vccd1 vccd1 _14935_/B sky130_fd_sc_hd__nor2_2
X_10049_ _10044_/A _10047_/X _10048_/X _10010_/A vssd1 vssd1 vccd1 vccd1 _10053_/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_209_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18694_ _18732_/CLK _18694_/D vssd1 vssd1 vccd1 vccd1 _18694_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_76_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17645_ _18184_/Q vssd1 vssd1 vccd1 vccd1 _17645_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_75_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14857_ _18303_/Q _14861_/B _14856_/X _14839_/X vssd1 vssd1 vccd1 vccd1 _18303_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_223_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13808_ _18393_/Q _13785_/A _13766_/A _18375_/Q vssd1 vssd1 vccd1 vccd1 _13808_/X
+ sky130_fd_sc_hd__a22o_1
X_14788_ _14814_/A _14788_/B vssd1 vssd1 vccd1 vccd1 _14788_/Y sky130_fd_sc_hd__nand2_1
X_17576_ _17602_/A _17674_/A vssd1 vssd1 vccd1 vccd1 _17576_/Y sky130_fd_sc_hd__nor2_2
XFILLER_91_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_220_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_205_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16527_ _16672_/A _16652_/C vssd1 vssd1 vccd1 vccd1 _16538_/B sky130_fd_sc_hd__nor2_1
X_13739_ _13781_/A vssd1 vssd1 vccd1 vccd1 _13739_/X sky130_fd_sc_hd__buf_8
XFILLER_91_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_220_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_220_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_220_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16458_ _18721_/Q _18685_/Q _16470_/S vssd1 vssd1 vccd1 vccd1 _16458_/X sky130_fd_sc_hd__mux2_1
XFILLER_108_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15409_ _16922_/A vssd1 vssd1 vccd1 vccd1 _16007_/B sky130_fd_sc_hd__buf_2
X_16389_ _16389_/A _16392_/B vssd1 vssd1 vccd1 vccd1 _16389_/Y sky130_fd_sc_hd__nand2_1
XFILLER_191_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19177_ _19177_/A _09009_/Y vssd1 vssd1 vccd1 vccd1 io_out[15] sky130_fd_sc_hd__ebufn_8
XFILLER_145_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18128_ _19027_/CLK _18128_/D vssd1 vssd1 vccd1 vccd1 _18128_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_172_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_117_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18059_ _18069_/CLK _18059_/D vssd1 vssd1 vccd1 vccd1 _18059_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_132_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09901_ _09901_/A _09907_/A vssd1 vssd1 vccd1 vccd1 _09910_/B sky130_fd_sc_hd__nand2_1
XFILLER_28_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_141_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09832_ _12112_/B _12112_/C vssd1 vssd1 vccd1 vccd1 _09833_/B sky130_fd_sc_hd__xor2_1
XFILLER_8_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09763_ _17784_/Q vssd1 vssd1 vccd1 vccd1 _09792_/A sky130_fd_sc_hd__clkinv_2
XFILLER_39_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_227_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09694_ _09694_/A vssd1 vssd1 vccd1 vccd1 _09711_/A sky130_fd_sc_hd__buf_4
XFILLER_227_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_230_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_212_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_230_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_223_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_211_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_136_wb_clk_i clkbuf_5_27_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18346_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_228_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_1288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_194_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09128_ _18827_/Q _18826_/Q _18825_/Q vssd1 vssd1 vccd1 vccd1 _09131_/B sky130_fd_sc_hd__or3_4
XFILLER_157_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_191_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09059_ _11018_/A vssd1 vssd1 vccd1 vccd1 _09059_/Y sky130_fd_sc_hd__inv_2
XFILLER_194_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_1340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12070_ _12070_/A _12070_/B vssd1 vssd1 vccd1 vccd1 _12070_/Y sky130_fd_sc_hd__nor2_1
XFILLER_2_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11021_ _13344_/A vssd1 vssd1 vccd1 vccd1 _11021_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_77_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_1316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15760_ _15821_/A vssd1 vssd1 vccd1 vccd1 _15892_/B sky130_fd_sc_hd__buf_2
XTAP_4144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12972_ _12972_/A vssd1 vssd1 vccd1 vccd1 _12972_/X sky130_fd_sc_hd__buf_4
XFILLER_218_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14711_ _14734_/A _15150_/B _14757_/C vssd1 vssd1 vccd1 vccd1 _14711_/X sky130_fd_sc_hd__or3_1
XFILLER_46_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11923_ _13509_/B vssd1 vssd1 vccd1 vccd1 _12126_/B sky130_fd_sc_hd__clkbuf_2
X_15691_ _15691_/A _15694_/B vssd1 vssd1 vccd1 vccd1 _15691_/Y sky130_fd_sc_hd__nand2_1
XFILLER_206_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14642_ _14665_/A _14665_/B _15233_/B vssd1 vssd1 vccd1 vccd1 _14642_/X sky130_fd_sc_hd__or3_1
XTAP_3498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17430_ _17543_/S vssd1 vssd1 vccd1 vccd1 _17447_/S sky130_fd_sc_hd__clkbuf_2
XTAP_2753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11854_ _17517_/A vssd1 vssd1 vccd1 vccd1 _14185_/A sky130_fd_sc_hd__buf_6
XTAP_2764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10805_ _10805_/A _10805_/B _10805_/C vssd1 vssd1 vccd1 vccd1 _10805_/X sky130_fd_sc_hd__and3_1
X_14573_ _18238_/Q _14574_/B _14572_/Y _14561_/X vssd1 vssd1 vccd1 vccd1 _18238_/D
+ sky130_fd_sc_hd__o211a_1
X_17361_ _17400_/A vssd1 vssd1 vccd1 vccd1 _17361_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_198_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11785_ _13446_/A _13429_/A vssd1 vssd1 vccd1 vccd1 _11786_/A sky130_fd_sc_hd__nand2_1
XFILLER_60_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_198_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16312_ _18685_/Q _18649_/Q _16324_/S vssd1 vssd1 vccd1 vccd1 _16312_/X sky130_fd_sc_hd__mux2_1
X_13524_ _13524_/A vssd1 vssd1 vccd1 vccd1 _13525_/A sky130_fd_sc_hd__buf_4
XFILLER_207_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10736_ _09093_/C _09098_/B _10882_/S vssd1 vssd1 vccd1 vccd1 _10736_/X sky130_fd_sc_hd__mux2_1
X_17292_ _17291_/B _17289_/X _17291_/Y _17283_/X vssd1 vssd1 vccd1 vccd1 _18884_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_198_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16243_ _16268_/A _16243_/B vssd1 vssd1 vccd1 vccd1 _16243_/Y sky130_fd_sc_hd__nand2_1
X_19031_ _19031_/CLK _19031_/D vssd1 vssd1 vccd1 vccd1 _19031_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_186_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13455_ _13455_/A _13455_/B _13455_/C vssd1 vssd1 vccd1 vccd1 _13456_/C sky130_fd_sc_hd__nor3_1
XFILLER_40_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10667_ _10667_/A vssd1 vssd1 vccd1 vccd1 _10671_/B sky130_fd_sc_hd__buf_2
X_12406_ _12406_/A _12406_/B _12406_/C vssd1 vssd1 vccd1 vccd1 _12407_/C sky130_fd_sc_hd__or3_1
X_16174_ _18653_/Q _18617_/Q _16192_/S vssd1 vssd1 vccd1 vccd1 _16174_/X sky130_fd_sc_hd__mux2_1
XFILLER_51_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13386_ _17972_/Q _17971_/Q vssd1 vssd1 vccd1 vccd1 _13386_/Y sky130_fd_sc_hd__nor2_1
XFILLER_103_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10598_ _10598_/A _10598_/B vssd1 vssd1 vccd1 vccd1 _10598_/X sky130_fd_sc_hd__or2_1
X_15125_ _15125_/A vssd1 vssd1 vccd1 vccd1 _15141_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_127_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_217_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12337_ _12328_/B _12336_/X _12337_/S vssd1 vssd1 vccd1 vccd1 _12338_/B sky130_fd_sc_hd__mux2_1
XFILLER_126_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_181_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15056_ _15105_/A vssd1 vssd1 vccd1 vccd1 _15081_/S sky130_fd_sc_hd__clkbuf_2
X_12268_ _12147_/X _11569_/B _12266_/X _12267_/X vssd1 vssd1 vccd1 vccd1 _17866_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_123_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14007_ _12022_/C _13999_/X _14006_/X _12027_/D vssd1 vssd1 vccd1 vccd1 _14007_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_218_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11219_ _17816_/Q _11215_/B _11218_/X vssd1 vssd1 vccd1 vccd1 _11220_/B sky130_fd_sc_hd__o21ai_1
XFILLER_214_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12199_ _12493_/B _12358_/B vssd1 vssd1 vccd1 vccd1 _12205_/A sky130_fd_sc_hd__nor2_1
XFILLER_150_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18815_ _18826_/CLK _18815_/D vssd1 vssd1 vccd1 vccd1 _18815_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_68_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18746_ _18752_/CLK _18746_/D vssd1 vssd1 vccd1 vccd1 _18746_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_5390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15958_ _17228_/A vssd1 vssd1 vccd1 vccd1 _16216_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_3_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_224_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14909_ _18352_/Q _18316_/Q _14934_/S vssd1 vssd1 vccd1 vccd1 _14909_/X sky130_fd_sc_hd__mux2_1
XFILLER_3_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18677_ _18677_/CLK _18677_/D vssd1 vssd1 vccd1 vccd1 _18677_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_64_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15889_ _15889_/A vssd1 vssd1 vccd1 vccd1 _15942_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_36_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_1277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_224_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17628_ _17567_/X _17623_/Y _17603_/X _17624_/Y _18970_/Q vssd1 vssd1 vccd1 vccd1
+ _17629_/B sky130_fd_sc_hd__a32o_1
XFILLER_23_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_196_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_225_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17559_ _14360_/X _16975_/A _17547_/X _17558_/X _17556_/X vssd1 vssd1 vccd1 vccd1
+ _18953_/D sky130_fd_sc_hd__o311a_1
XFILLER_32_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_221_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19229_ _19229_/A _08941_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[29] sky130_fd_sc_hd__ebufn_8
XFILLER_176_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_145_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_207_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09815_ _09813_/A _09795_/Y _09797_/Y vssd1 vssd1 vccd1 vccd1 _09818_/A sky130_fd_sc_hd__a21o_1
XFILLER_100_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19054__25 vssd1 vssd1 vccd1 vccd1 _19054__25/HI _19148_/A sky130_fd_sc_hd__conb_1
XFILLER_115_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_189_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_228_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09746_ _09752_/A _09746_/B vssd1 vssd1 vccd1 vccd1 _09748_/C sky130_fd_sc_hd__xnor2_1
XFILLER_27_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_227_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09677_ _18236_/Q _18235_/Q _18234_/Q vssd1 vssd1 vccd1 vccd1 _09677_/X sky130_fd_sc_hd__or3_4
XTAP_2016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_161_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11570_ _11570_/A _11570_/B vssd1 vssd1 vccd1 vccd1 _11570_/X sky130_fd_sc_hd__or2_1
XFILLER_139_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_210_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10521_ _10521_/A vssd1 vssd1 vccd1 vccd1 _10522_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_122_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_1361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13240_ _13244_/A _18075_/Q vssd1 vssd1 vccd1 vccd1 _13241_/A sky130_fd_sc_hd__and2_1
XFILLER_202_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10452_ _10450_/X _10451_/X _10496_/A vssd1 vssd1 vccd1 vccd1 _10452_/X sky130_fd_sc_hd__mux2_2
X_13171_ _13175_/A _18044_/Q vssd1 vssd1 vccd1 vccd1 _13172_/A sky130_fd_sc_hd__and2_1
XFILLER_163_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10383_ _09309_/D _10316_/S _10382_/X _09937_/X vssd1 vssd1 vccd1 vccd1 _10383_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_123_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_33_wb_clk_i clkbuf_5_18_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18245_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_11_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12122_ _12122_/A _13420_/A vssd1 vssd1 vccd1 vccd1 _12127_/B sky130_fd_sc_hd__nor2_1
XFILLER_184_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16930_ _16957_/A _16930_/B vssd1 vssd1 vccd1 vccd1 _16930_/Y sky130_fd_sc_hd__nand2_1
XFILLER_123_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12053_ _12053_/A _12053_/B _13710_/A vssd1 vssd1 vccd1 vccd1 _12054_/D sky130_fd_sc_hd__and3_1
XFILLER_105_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_1271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11004_ _11232_/A _11232_/B _11001_/C _11003_/X vssd1 vssd1 vccd1 vccd1 _19173_/A
+ sky130_fd_sc_hd__o31ai_4
XFILLER_89_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16861_ _16860_/B _16859_/X _16860_/Y _16848_/X vssd1 vssd1 vccd1 vccd1 _18782_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_78_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18600_ _18635_/CLK _18600_/D vssd1 vssd1 vccd1 vccd1 _18600_/Q sky130_fd_sc_hd__dfxtp_4
X_15812_ _15818_/B _15809_/X _15811_/X _15803_/X vssd1 vssd1 vccd1 vccd1 _18531_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_77_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16792_ _16815_/A _16792_/B vssd1 vssd1 vccd1 vccd1 _16792_/Y sky130_fd_sc_hd__nand2_1
XFILLER_92_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_206_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18531_ _18533_/CLK _18531_/D vssd1 vssd1 vccd1 vccd1 _18531_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_219_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15743_ _15754_/A _15743_/B vssd1 vssd1 vccd1 vccd1 _15743_/Y sky130_fd_sc_hd__nand2_1
XTAP_3240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12955_ _12955_/A vssd1 vssd1 vccd1 vccd1 _12955_/X sky130_fd_sc_hd__clkbuf_2
XTAP_3251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11906_ _12142_/A vssd1 vssd1 vccd1 vccd1 _12141_/A sky130_fd_sc_hd__inv_2
XFILLER_18_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18462_ _18485_/CLK _18462_/D vssd1 vssd1 vccd1 vccd1 _18462_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15674_ _15673_/B _15672_/X _15673_/Y _15662_/X vssd1 vssd1 vccd1 vccd1 _18497_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_206_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12886_ _17958_/Q _17959_/Q _12886_/C vssd1 vssd1 vccd1 vccd1 _12890_/B sky130_fd_sc_hd__and3_1
XTAP_2550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17413_ _17472_/A vssd1 vssd1 vccd1 vccd1 _17536_/B sky130_fd_sc_hd__buf_2
X_14625_ _14651_/A _15218_/A vssd1 vssd1 vccd1 vccd1 _14635_/B sky130_fd_sc_hd__nor2_1
X_11837_ _11484_/B _11836_/X _11488_/Y vssd1 vssd1 vccd1 vccd1 _11837_/X sky130_fd_sc_hd__o21a_1
XFILLER_33_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18393_ _18393_/CLK _18393_/D vssd1 vssd1 vccd1 vccd1 _18393_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_2594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14556_ _18234_/Q _14559_/B _14555_/X _14533_/X vssd1 vssd1 vccd1 vccd1 _18234_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_1893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17344_ _17464_/A vssd1 vssd1 vccd1 vccd1 _17392_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_198_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_158_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11768_ _11761_/A _11760_/B _11767_/A vssd1 vssd1 vccd1 vccd1 _11781_/B sky130_fd_sc_hd__a21oi_1
XFILLER_53_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13507_ _13507_/A vssd1 vssd1 vccd1 vccd1 _13508_/A sky130_fd_sc_hd__buf_6
XFILLER_159_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10719_ _10810_/S vssd1 vssd1 vccd1 vccd1 _10841_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_158_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14487_ _18218_/Q _14491_/B vssd1 vssd1 vccd1 vccd1 _14488_/A sky130_fd_sc_hd__and2_1
X_17275_ _17275_/A _17275_/B vssd1 vssd1 vccd1 vccd1 _17275_/Y sky130_fd_sc_hd__nand2_1
XFILLER_186_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11699_ _17852_/Q vssd1 vssd1 vccd1 vccd1 _11704_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_105_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_228_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_220_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19014_ _19029_/CLK _19014_/D vssd1 vssd1 vccd1 vccd1 _19014_/Q sky130_fd_sc_hd__dfxtp_1
X_16226_ _18627_/Q _16229_/B _16225_/X _16209_/X vssd1 vssd1 vccd1 vccd1 _18627_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_146_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13438_ _13438_/A _13438_/B _13438_/C vssd1 vssd1 vccd1 vccd1 _13439_/B sky130_fd_sc_hd__or3_1
XFILLER_220_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16157_ _16199_/A _16160_/B vssd1 vssd1 vccd1 vccd1 _16157_/Y sky130_fd_sc_hd__nand2_1
XFILLER_127_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13369_ _10123_/A _13337_/X _13368_/Y vssd1 vssd1 vccd1 vccd1 _13370_/C sky130_fd_sc_hd__a21o_1
XFILLER_138_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15108_ _15107_/B _15106_/X _15107_/Y _15103_/X vssd1 vssd1 vccd1 vccd1 _18365_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_138_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16088_ _16839_/A vssd1 vssd1 vccd1 vccd1 _16692_/B sky130_fd_sc_hd__buf_4
XFILLER_103_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15039_ _15038_/B _15037_/X _15038_/Y _15026_/X vssd1 vssd1 vccd1 vccd1 _18347_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_218_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_1311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_1243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_1306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09600_ _09600_/A _09600_/B _09600_/C vssd1 vssd1 vccd1 vccd1 _09601_/B sky130_fd_sc_hd__and3_1
XFILLER_96_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_216_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09531_ _18125_/Q _09531_/B vssd1 vssd1 vccd1 vccd1 _09568_/A sky130_fd_sc_hd__xor2_4
XFILLER_209_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18729_ _18738_/CLK _18729_/D vssd1 vssd1 vccd1 vccd1 _18729_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_64_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09462_ _09462_/A vssd1 vssd1 vccd1 vccd1 _18132_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_19_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_149_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09393_ _18374_/Q _18373_/Q _18372_/Q vssd1 vssd1 vccd1 vccd1 _09397_/A sky130_fd_sc_hd__or3_4
XFILLER_24_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_225_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_4_1_0_wb_clk_i clkbuf_4_1_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_5_3_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_156_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_219_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_219_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09729_ _17784_/Q vssd1 vssd1 vccd1 vccd1 _09802_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_210_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12740_ _19008_/Q _19007_/Q _19010_/Q _19009_/Q vssd1 vssd1 vccd1 vccd1 _12742_/B
+ sky130_fd_sc_hd__and4_1
XTAP_1101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_231_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12671_ _12671_/A vssd1 vssd1 vccd1 vccd1 _12672_/B sky130_fd_sc_hd__inv_2
XTAP_1156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_230_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14410_ _14404_/A _14409_/B _14423_/A vssd1 vssd1 vccd1 vccd1 _14410_/X sky130_fd_sc_hd__a21o_1
XFILLER_208_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11622_ _11622_/A vssd1 vssd1 vccd1 vccd1 _11689_/A sky130_fd_sc_hd__clkbuf_2
X_15390_ _15445_/A _15390_/B vssd1 vssd1 vccd1 vccd1 _15390_/Y sky130_fd_sc_hd__nand2_1
XTAP_1189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_230_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14341_ _14275_/X _14337_/X _14339_/X _14340_/X vssd1 vssd1 vccd1 vccd1 _18179_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_169_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11553_ _11562_/A _17865_/Q vssd1 vssd1 vccd1 vccd1 _11553_/Y sky130_fd_sc_hd__nor2_1
XFILLER_195_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10504_ _09143_/D _09148_/A _10550_/S vssd1 vssd1 vccd1 vccd1 _10504_/X sky130_fd_sc_hd__mux2_1
X_17060_ _17078_/A vssd1 vssd1 vccd1 vccd1 _17074_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_7_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14272_ _14272_/A _14272_/B _14283_/A vssd1 vssd1 vccd1 vccd1 _14272_/X sky130_fd_sc_hd__and3_2
XFILLER_156_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11484_ _11484_/A _11484_/B vssd1 vssd1 vccd1 vccd1 _11484_/X sky130_fd_sc_hd__and2_1
X_16011_ _16212_/A vssd1 vssd1 vccd1 vccd1 _16062_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_7_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13223_ _13223_/A vssd1 vssd1 vccd1 vccd1 _18066_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_13_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10435_ _10427_/X _10434_/X _10918_/S vssd1 vssd1 vccd1 vccd1 _10436_/C sky130_fd_sc_hd__mux2_1
XFILLER_100_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_1333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13154_ _16891_/A vssd1 vssd1 vccd1 vccd1 _13199_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_3_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10366_ _10403_/A _10366_/B vssd1 vssd1 vccd1 vccd1 _10366_/X sky130_fd_sc_hd__and2b_1
XFILLER_152_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12105_ _12056_/Y _12069_/X _12085_/Y _12088_/X _12104_/X vssd1 vssd1 vccd1 vccd1
+ _12105_/X sky130_fd_sc_hd__o41a_1
XFILLER_97_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13085_ _13085_/A _14480_/B vssd1 vssd1 vccd1 vccd1 _13086_/A sky130_fd_sc_hd__and2_1
X_17962_ _17965_/CLK _17962_/D vssd1 vssd1 vccd1 vccd1 _17962_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_88_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10297_ _10305_/S _10290_/X _10296_/X _09895_/X vssd1 vssd1 vccd1 vccd1 _10312_/A
+ sky130_fd_sc_hd__o211a_1
X_16913_ _16954_/A _16916_/B vssd1 vssd1 vccd1 vccd1 _16913_/Y sky130_fd_sc_hd__nand2_1
X_12036_ _17803_/Q _12036_/B vssd1 vssd1 vccd1 vccd1 _12037_/B sky130_fd_sc_hd__nand2_1
XFILLER_78_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17893_ _17895_/CLK _17893_/D vssd1 vssd1 vccd1 vccd1 _17893_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_215_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16844_ _16847_/B _16842_/X _16843_/Y _16825_/X vssd1 vssd1 vccd1 vccd1 _18778_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_38_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16775_ _18799_/Q _18763_/Q _16784_/S vssd1 vssd1 vccd1 vccd1 _16775_/X sky130_fd_sc_hd__mux2_1
XFILLER_4_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13987_ _18397_/Q _13583_/A _13489_/A _18388_/Q vssd1 vssd1 vccd1 vccd1 _13987_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_34_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_230_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18514_ _18553_/CLK _18514_/D vssd1 vssd1 vccd1 vccd1 _18514_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15726_ _18547_/Q _18511_/Q _15733_/S vssd1 vssd1 vccd1 vccd1 _15726_/X sky130_fd_sc_hd__mux2_1
XFILLER_19_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12938_ _11025_/B _12933_/A _12764_/X vssd1 vssd1 vccd1 vccd1 _12939_/B sky130_fd_sc_hd__o21ai_1
XFILLER_59_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_222_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_146_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_209_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18445_ _18448_/CLK _18445_/D vssd1 vssd1 vccd1 vccd1 _18445_/Q sky130_fd_sc_hd__dfxtp_1
X_15657_ _18529_/Q _18493_/Q _15665_/S vssd1 vssd1 vccd1 vccd1 _15657_/X sky130_fd_sc_hd__mux2_1
XFILLER_181_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12869_ _12869_/A vssd1 vssd1 vccd1 vccd1 _12871_/B sky130_fd_sc_hd__inv_2
XTAP_2391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14608_ _14687_/A vssd1 vssd1 vccd1 vccd1 _14608_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_222_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18376_ _18408_/CLK _18376_/D vssd1 vssd1 vccd1 vccd1 _18376_/Q sky130_fd_sc_hd__dfxtp_1
X_15588_ _15594_/B _15586_/X _15587_/X _15575_/X vssd1 vssd1 vccd1 vccd1 _18477_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_159_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_175_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17327_ _17336_/A _17327_/B vssd1 vssd1 vccd1 vccd1 _17327_/Y sky130_fd_sc_hd__nand2_1
X_14539_ _14604_/A _14545_/B vssd1 vssd1 vccd1 vccd1 _14539_/Y sky130_fd_sc_hd__nand2_1
XFILLER_175_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_179_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17258_ _18913_/Q _18877_/Q _17262_/S vssd1 vssd1 vccd1 vccd1 _17258_/X sky130_fd_sc_hd__mux2_1
XFILLER_105_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16209_ _16252_/A vssd1 vssd1 vccd1 vccd1 _16209_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_179_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17189_ _17213_/A _17189_/B vssd1 vssd1 vccd1 vccd1 _17189_/Y sky130_fd_sc_hd__nand2_1
XFILLER_115_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_1302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08962_ _08966_/A vssd1 vssd1 vccd1 vccd1 _08962_/Y sky130_fd_sc_hd__inv_2
XFILLER_130_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_229_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_112_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_216_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09514_ _18227_/Q _14372_/B vssd1 vssd1 vccd1 vccd1 _14510_/B sky130_fd_sc_hd__or2_1
XFILLER_140_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_231_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_225_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09445_ _09188_/A _09187_/Y _09430_/D vssd1 vssd1 vccd1 vccd1 _09445_/Y sky130_fd_sc_hd__o21ai_1
XPHY_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_227_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_212_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09376_ _09376_/A _09376_/B _09376_/C _09376_/D vssd1 vssd1 vccd1 vccd1 _09387_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_197_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_200_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_221_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10220_ _10221_/B _10220_/B vssd1 vssd1 vccd1 vccd1 _10232_/B sky130_fd_sc_hd__xnor2_2
XFILLER_165_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10151_ _18119_/Q vssd1 vssd1 vccd1 vccd1 _13389_/A sky130_fd_sc_hd__clkbuf_2
XTAP_5901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10082_ _09287_/A _09287_/D _09282_/D _09282_/B _09703_/A _09709_/A vssd1 vssd1 vccd1
+ vccd1 _10082_/X sky130_fd_sc_hd__mux4_1
XTAP_5934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13910_ _18868_/Q _13529_/A _13725_/X _18844_/Q vssd1 vssd1 vccd1 vccd1 _13910_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_5978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14890_ _14935_/A _14890_/B vssd1 vssd1 vccd1 vccd1 _14890_/Y sky130_fd_sc_hd__nand2_1
XFILLER_134_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13841_ _13841_/A vssd1 vssd1 vccd1 vccd1 _13842_/A sky130_fd_sc_hd__buf_8
XFILLER_74_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16560_ _16562_/B _16557_/X _16558_/Y _16559_/X vssd1 vssd1 vccd1 vccd1 _18709_/D
+ sky130_fd_sc_hd__o211a_1
X_13772_ _13772_/A vssd1 vssd1 vccd1 vccd1 _13772_/X sky130_fd_sc_hd__buf_6
XFILLER_15_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_222_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10984_ _14187_/A vssd1 vssd1 vccd1 vccd1 _14317_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_204_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_215_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15511_ _15511_/A _15511_/B vssd1 vssd1 vccd1 vccd1 _15511_/Y sky130_fd_sc_hd__nand2_1
XFILLER_204_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12723_ _18001_/Q vssd1 vssd1 vccd1 vccd1 _12781_/B sky130_fd_sc_hd__inv_2
X_16491_ _16491_/A _16785_/B _16504_/C vssd1 vssd1 vccd1 vccd1 _16491_/X sky130_fd_sc_hd__or3_1
XFILLER_71_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18230_ _18230_/CLK _18230_/D vssd1 vssd1 vccd1 vccd1 _18230_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_70_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15442_ _15442_/A _15445_/B vssd1 vssd1 vccd1 vccd1 _15442_/Y sky130_fd_sc_hd__nand2_1
X_12654_ _12654_/A _12654_/B vssd1 vssd1 vccd1 vccd1 _12656_/A sky130_fd_sc_hd__nor2_1
XFILLER_128_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11605_ _17855_/Q vssd1 vssd1 vccd1 vccd1 _11624_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_156_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18161_ _19021_/CLK _18161_/D vssd1 vssd1 vccd1 vccd1 _18161_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_230_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15373_ _15373_/A _15375_/B vssd1 vssd1 vccd1 vccd1 _15373_/Y sky130_fd_sc_hd__nand2_1
XFILLER_156_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12585_ _17922_/Q _12569_/X _12589_/B _12584_/Y _12548_/X vssd1 vssd1 vccd1 vccd1
+ _17922_/D sky130_fd_sc_hd__a221o_1
XFILLER_196_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17112_ _17152_/A _17115_/B vssd1 vssd1 vccd1 vccd1 _17112_/Y sky130_fd_sc_hd__nand2_1
XFILLER_156_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11536_ _19031_/Q _11527_/Y _11528_/X _11535_/X vssd1 vssd1 vccd1 vccd1 _11536_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_11_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14324_ _14335_/B _18209_/Q vssd1 vssd1 vccd1 vccd1 _14325_/B sky130_fd_sc_hd__and2b_1
X_18092_ _18224_/CLK _18092_/D vssd1 vssd1 vccd1 vccd1 _18092_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_89_1338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_209_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17043_ _17088_/A _17046_/B vssd1 vssd1 vccd1 vccd1 _17043_/Y sky130_fd_sc_hd__nand2_1
X_14255_ _14202_/X _14253_/X _14254_/X _13334_/X vssd1 vssd1 vccd1 vccd1 _18171_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_143_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11467_ _11452_/A _11593_/A _11467_/C _11467_/D vssd1 vssd1 vccd1 vccd1 _11482_/B
+ sky130_fd_sc_hd__and4b_1
XFILLER_99_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13206_ _13208_/A _18060_/Q vssd1 vssd1 vccd1 vccd1 _13207_/A sky130_fd_sc_hd__and2_1
XFILLER_109_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10418_ _09209_/C _09214_/C _09219_/A _10795_/A _10236_/A _10413_/X vssd1 vssd1 vccd1
+ vccd1 _10419_/B sky130_fd_sc_hd__mux4_2
XFILLER_171_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14186_ _13412_/A _13412_/B _13418_/D _17941_/Q vssd1 vssd1 vccd1 vccd1 _14355_/C
+ sky130_fd_sc_hd__a211o_2
X_11398_ _11506_/B _11542_/B _13485_/A vssd1 vssd1 vccd1 vccd1 _11399_/A sky130_fd_sc_hd__o21a_1
XFILLER_48_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_180_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13137_ _13137_/A vssd1 vssd1 vccd1 vccd1 _18027_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_225_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10349_ _09119_/A _09109_/D _10349_/S vssd1 vssd1 vccd1 vccd1 _10349_/X sky130_fd_sc_hd__mux2_1
XTAP_715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18994_ _19000_/CLK _18994_/D vssd1 vssd1 vccd1 vccd1 _18994_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_97_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13068_ _18151_/Q _12927_/Y _12761_/X vssd1 vssd1 vccd1 vccd1 _13069_/S sky130_fd_sc_hd__o21a_1
X_17945_ _17959_/CLK _17945_/D vssd1 vssd1 vccd1 vccd1 _17945_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_215_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_227_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12019_ _12019_/A _12019_/B vssd1 vssd1 vccd1 vccd1 _12055_/D sky130_fd_sc_hd__or2_1
XFILLER_38_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17876_ _17879_/CLK _17876_/D vssd1 vssd1 vccd1 vccd1 _17876_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_17_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16827_ _18811_/Q _18775_/Q _16842_/S vssd1 vssd1 vccd1 vccd1 _16827_/X sky130_fd_sc_hd__mux2_1
XFILLER_54_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16758_ _18795_/Q _18759_/Q _16762_/S vssd1 vssd1 vccd1 vccd1 _16758_/X sky130_fd_sc_hd__mux2_1
XFILLER_81_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19037__8 vssd1 vssd1 vccd1 vccd1 _19037__8/HI _19131_/A sky130_fd_sc_hd__conb_1
XFILLER_34_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15709_ _15708_/B _15706_/X _15708_/Y _15700_/X vssd1 vssd1 vccd1 vccd1 _18506_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_185_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16689_ _16689_/A _16745_/B vssd1 vssd1 vccd1 vccd1 _16699_/B sky130_fd_sc_hd__nor2_2
XFILLER_224_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09230_ _18920_/Q _18919_/Q _18918_/Q vssd1 vssd1 vccd1 vccd1 _09232_/C sky130_fd_sc_hd__or3_4
X_18428_ _18434_/CLK _18428_/D vssd1 vssd1 vccd1 vccd1 _18428_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_21_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_222_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_181_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_1178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_222_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09161_ _18641_/Q _18640_/Q _18639_/Q vssd1 vssd1 vccd1 vccd1 _09165_/A sky130_fd_sc_hd__or3_4
XFILLER_148_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18359_ _18387_/CLK _18359_/D vssd1 vssd1 vccd1 vccd1 _18359_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_187_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_222_1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09092_ _18806_/Q _18805_/Q _18804_/Q vssd1 vssd1 vccd1 vccd1 _09093_/D sky130_fd_sc_hd__or3_4
XFILLER_120_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_175_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_1274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09994_ _10046_/A vssd1 vssd1 vccd1 vccd1 _09995_/A sky130_fd_sc_hd__buf_6
XFILLER_192_1176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08945_ _08948_/A vssd1 vssd1 vccd1 vccd1 _08945_/Y sky130_fd_sc_hd__inv_2
XFILLER_131_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_231_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_213_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_197_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_213_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09428_ _09450_/A _09420_/X _09427_/Y _09421_/Y _09221_/B vssd1 vssd1 vccd1 vccd1
+ _09428_/X sky130_fd_sc_hd__o311a_2
XFILLER_13_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_125_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_212_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_212_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09359_ _18290_/Q _18289_/Q _18288_/Q vssd1 vssd1 vccd1 vccd1 _09360_/D sky130_fd_sc_hd__or3_4
XFILLER_166_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12370_ _12370_/A vssd1 vssd1 vccd1 vccd1 _17893_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_121_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_165_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11321_ _11345_/A vssd1 vssd1 vccd1 vccd1 _11323_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_193_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_197_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_181_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14040_ _18335_/Q _13837_/A _14038_/X _14039_/X vssd1 vssd1 vccd1 vccd1 _14040_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_158_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11252_ _11788_/A _11735_/B _11455_/C vssd1 vssd1 vccd1 vccd1 _11396_/B sky130_fd_sc_hd__a21o_2
Xclkbuf_5_10_0_wb_clk_i clkbuf_4_5_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_5_10_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_141_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10203_ _18120_/Q vssd1 vssd1 vccd1 vccd1 _10206_/A sky130_fd_sc_hd__inv_2
XFILLER_45_1208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11183_ _11183_/A vssd1 vssd1 vccd1 vccd1 _17807_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_69_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_106_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10134_ _18127_/Q vssd1 vssd1 vccd1 vccd1 _10141_/A sky130_fd_sc_hd__inv_2
XFILLER_0_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15991_ _16003_/A _15991_/B vssd1 vssd1 vccd1 vccd1 _15991_/Y sky130_fd_sc_hd__nand2_1
XTAP_5731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17730_ _17734_/A _19010_/Q vssd1 vssd1 vccd1 vccd1 _17731_/A sky130_fd_sc_hd__and2_1
XFILLER_0_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14942_ _14949_/B _14939_/X _14940_/X _14941_/X vssd1 vssd1 vccd1 vccd1 _18324_/D
+ sky130_fd_sc_hd__o211a_1
X_10065_ _10065_/A _10065_/B _10065_/C vssd1 vssd1 vccd1 vccd1 _10065_/X sky130_fd_sc_hd__and3_1
XTAP_5764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17661_ _17661_/A vssd1 vssd1 vccd1 vccd1 _17736_/A sky130_fd_sc_hd__buf_4
X_14873_ _14875_/B _14871_/X _14872_/Y _14859_/X vssd1 vssd1 vccd1 vccd1 _18307_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_91_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_1290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16612_ _16611_/B _16610_/X _16611_/Y _16600_/X vssd1 vssd1 vccd1 vccd1 _18722_/D
+ sky130_fd_sc_hd__o211a_1
X_13824_ _18585_/Q _13657_/A _13822_/X _13823_/X vssd1 vssd1 vccd1 vccd1 _13824_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_75_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_1274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17592_ _17590_/Y _17552_/A _17591_/X vssd1 vssd1 vccd1 vccd1 _17592_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_90_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_105 _13877_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINSDIODE2_116 _16839_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINSDIODE2_127 _15279_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_138 _15440_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16543_ _18741_/Q _18705_/Q _16546_/S vssd1 vssd1 vccd1 vccd1 _16543_/X sky130_fd_sc_hd__mux2_1
XFILLER_182_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13755_ _18789_/Q _13522_/A _13753_/X _13754_/X vssd1 vssd1 vccd1 vccd1 _13755_/X
+ sky130_fd_sc_hd__a211o_1
X_10967_ _10938_/Y _10939_/X _10965_/Y _10966_/Y vssd1 vssd1 vccd1 vccd1 _13411_/D
+ sky130_fd_sc_hd__o22ai_2
XINSDIODE2_149 _18958_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12706_ _12707_/B _12707_/C _12707_/A vssd1 vssd1 vccd1 vccd1 _12708_/B sky130_fd_sc_hd__o21a_1
X_16474_ _18725_/Q _18689_/Q _16490_/S vssd1 vssd1 vccd1 vccd1 _16474_/X sky130_fd_sc_hd__mux2_1
XFILLER_231_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13686_ _18624_/Q _13758_/A _13697_/A _18615_/Q vssd1 vssd1 vccd1 vccd1 _13686_/X
+ sky130_fd_sc_hd__a22o_1
X_10898_ _09413_/D _09418_/C _09418_/A _09408_/D _10429_/X _10484_/X vssd1 vssd1 vccd1
+ vccd1 _10899_/B sky130_fd_sc_hd__mux4_2
XFILLER_188_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18213_ _18213_/CLK _18213_/D vssd1 vssd1 vccd1 vccd1 _18213_/Q sky130_fd_sc_hd__dfxtp_1
X_15425_ _18475_/Q _18439_/Q _15435_/S vssd1 vssd1 vccd1 vccd1 _15425_/X sky130_fd_sc_hd__mux2_1
XFILLER_54_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19193_ _19193_/A _08994_/Y vssd1 vssd1 vccd1 vccd1 io_out[31] sky130_fd_sc_hd__ebufn_8
X_12637_ _17931_/Q _12637_/B vssd1 vssd1 vccd1 vccd1 _12638_/B sky130_fd_sc_hd__and2_1
XFILLER_19_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18144_ _18144_/CLK _18144_/D vssd1 vssd1 vccd1 vccd1 _18144_/Q sky130_fd_sc_hd__dfxtp_1
X_15356_ _18459_/Q _18423_/Q _15356_/S vssd1 vssd1 vccd1 vccd1 _15356_/X sky130_fd_sc_hd__mux2_1
XFILLER_15_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12568_ _12570_/B _12529_/X _12566_/Y _12567_/X _11896_/X vssd1 vssd1 vccd1 vccd1
+ _17920_/D sky130_fd_sc_hd__o221ai_1
XFILLER_106_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11519_ _11522_/A _11530_/B _11645_/A _12285_/B _12287_/A vssd1 vssd1 vccd1 vccd1
+ _11519_/X sky130_fd_sc_hd__o221a_1
X_14307_ _14307_/A _14307_/B vssd1 vssd1 vccd1 vccd1 _14307_/Y sky130_fd_sc_hd__nor2_1
XFILLER_89_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18075_ _18085_/CLK _18075_/D vssd1 vssd1 vccd1 vccd1 _18075_/Q sky130_fd_sc_hd__dfxtp_1
X_15287_ _15286_/B _15285_/X _15286_/Y _15283_/X vssd1 vssd1 vccd1 vccd1 _18410_/D
+ sky130_fd_sc_hd__o211a_1
X_12499_ _17908_/Q _17907_/Q _12499_/C _12499_/D vssd1 vssd1 vccd1 vccd1 _12499_/X
+ sky130_fd_sc_hd__and4_1
XFILLER_7_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17026_ _18855_/Q _18819_/Q _17026_/S vssd1 vssd1 vccd1 vccd1 _17026_/X sky130_fd_sc_hd__mux2_1
XFILLER_176_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14238_ _14317_/A _10948_/S _10852_/X _14237_/X vssd1 vssd1 vccd1 vccd1 _14238_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_172_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14169_ _18614_/Q _13856_/X _13493_/X _18605_/Q _14168_/X vssd1 vssd1 vccd1 vccd1
+ _14169_/X sky130_fd_sc_hd__a221o_1
XFILLER_124_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_112_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18977_ _18977_/CLK _18977_/D vssd1 vssd1 vccd1 vccd1 _18977_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_230_1302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17928_ _17931_/CLK _17928_/D vssd1 vssd1 vccd1 vccd1 _17928_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_227_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_230_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_227_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17859_ _17891_/CLK _17859_/D vssd1 vssd1 vccd1 vccd1 _17859_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_67_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_226_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_226_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_228_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_201_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_224_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_228_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09213_ _18689_/Q _18688_/Q _18687_/Q vssd1 vssd1 vccd1 vccd1 _09214_/D sky130_fd_sc_hd__or3_4
XFILLER_179_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_210_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09144_ _18734_/Q _18733_/Q _18732_/Q vssd1 vssd1 vccd1 vccd1 _09148_/A sky130_fd_sc_hd__or3_4
XFILLER_147_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09075_ _09083_/A _09081_/B _17830_/Q vssd1 vssd1 vccd1 vccd1 _09076_/A sky130_fd_sc_hd__and3_1
XFILLER_108_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_135_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09977_ _14260_/B _09968_/X _09975_/X _10605_/B vssd1 vssd1 vccd1 vccd1 _09977_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_5027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08928_ input1/X vssd1 vssd1 vccd1 vccd1 _09053_/A sky130_fd_sc_hd__buf_4
XTAP_4326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_58_wb_clk_i _18759_/CLK vssd1 vssd1 vccd1 vccd1 _18743_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_3658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11870_ _11868_/X _11869_/Y _11867_/A vssd1 vssd1 vccd1 vccd1 _11870_/Y sky130_fd_sc_hd__a21oi_4
XTAP_3669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10821_ _13009_/A _10821_/B vssd1 vssd1 vccd1 vccd1 _14330_/A sky130_fd_sc_hd__xnor2_4
XTAP_2957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13540_ _18687_/Q _13576_/A _13539_/X _18663_/Q vssd1 vssd1 vccd1 vccd1 _13540_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_13_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10752_ _13007_/A _10843_/B _10752_/C vssd1 vssd1 vccd1 vccd1 _10752_/X sky130_fd_sc_hd__and3_1
XFILLER_207_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13471_ _13480_/A _13471_/B vssd1 vssd1 vccd1 vccd1 _18158_/D sky130_fd_sc_hd__nor2_1
XFILLER_40_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10683_ _10809_/A vssd1 vssd1 vccd1 vccd1 _10824_/A sky130_fd_sc_hd__buf_4
XFILLER_90_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15210_ _15527_/A _15279_/C vssd1 vssd1 vccd1 vccd1 _15216_/B sky130_fd_sc_hd__nor2_2
XFILLER_185_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12422_ _12412_/A _12413_/X _12439_/A _12420_/X vssd1 vssd1 vccd1 vccd1 _12430_/B
+ sky130_fd_sc_hd__o211ai_2
XFILLER_71_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16190_ _16945_/A vssd1 vssd1 vccd1 vccd1 _16783_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_51_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_200_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15141_ _18410_/Q _18374_/Q _15141_/S vssd1 vssd1 vccd1 vccd1 _15141_/X sky130_fd_sc_hd__mux2_1
X_12353_ _12353_/A vssd1 vssd1 vccd1 vccd1 _12353_/Y sky130_fd_sc_hd__inv_2
XFILLER_51_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_142_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11304_ _17804_/Q _11501_/C _13509_/A vssd1 vssd1 vccd1 vccd1 _11488_/A sky130_fd_sc_hd__or3b_1
X_15072_ _15118_/A _15072_/B vssd1 vssd1 vccd1 vccd1 _15072_/Y sky130_fd_sc_hd__nand2_1
XFILLER_153_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12284_ _12304_/A _12304_/B vssd1 vssd1 vccd1 vccd1 _12284_/X sky130_fd_sc_hd__and2b_1
XFILLER_153_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14023_ _18860_/Q _13834_/X _14021_/X _14022_/X vssd1 vssd1 vccd1 vccd1 _14023_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_4_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18900_ _18902_/CLK _18900_/D vssd1 vssd1 vccd1 vccd1 _18900_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_136_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11235_ _11001_/C _11234_/A _11221_/X vssd1 vssd1 vccd1 vccd1 _11235_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_106_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18831_ _18849_/CLK _18831_/D vssd1 vssd1 vccd1 vccd1 _18831_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_150_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11166_ _17814_/Q vssd1 vssd1 vccd1 vccd1 _11209_/A sky130_fd_sc_hd__inv_2
XFILLER_96_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10117_ _10142_/A _10142_/B vssd1 vssd1 vccd1 vccd1 _10118_/B sky130_fd_sc_hd__xor2_1
Xclkbuf_4_14_0_wb_clk_i clkbuf_3_7_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_5_29_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_2
X_18762_ _18765_/CLK _18762_/D vssd1 vssd1 vccd1 vccd1 _18762_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_96_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15974_ _16287_/A _16043_/C vssd1 vssd1 vccd1 vccd1 _15980_/B sky130_fd_sc_hd__nor2_2
XTAP_5550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11097_ _17794_/Q vssd1 vssd1 vccd1 vccd1 _11281_/A sky130_fd_sc_hd__clkbuf_2
XTAP_5561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_222_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17713_ _17713_/A vssd1 vssd1 vccd1 vccd1 _19001_/D sky130_fd_sc_hd__clkbuf_1
XTAP_5583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10048_ _09186_/B _09176_/B _09181_/C _09186_/C _10036_/X _10956_/B vssd1 vssd1 vccd1
+ vccd1 _10048_/X sky130_fd_sc_hd__mux4_1
X_14925_ _18320_/Q _14924_/B _14924_/Y _14922_/X vssd1 vssd1 vccd1 vccd1 _18320_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_5594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18693_ _18693_/CLK _18693_/D vssd1 vssd1 vccd1 vccd1 _18693_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_48_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17644_ _17644_/A vssd1 vssd1 vccd1 vccd1 _18973_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14856_ _14856_/A _15150_/B _14906_/C vssd1 vssd1 vccd1 vccd1 _14856_/X sky130_fd_sc_hd__or3_1
XFILLER_1_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_223_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13807_ _18378_/Q _13677_/X _13764_/A _18402_/Q vssd1 vssd1 vccd1 vccd1 _13807_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_90_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17575_ _17575_/A vssd1 vssd1 vccd1 vccd1 _17575_/X sky130_fd_sc_hd__buf_2
X_14787_ _18323_/Q _18287_/Q _14787_/S vssd1 vssd1 vccd1 vccd1 _14787_/X sky130_fd_sc_hd__mux2_1
XFILLER_51_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11999_ _12041_/C _11999_/B _11999_/C vssd1 vssd1 vccd1 vccd1 _12006_/B sky130_fd_sc_hd__or3_1
XFILLER_95_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16526_ _18701_/Q _16525_/B _16525_/Y _16519_/X vssd1 vssd1 vccd1 vccd1 _18701_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_91_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13738_ _13738_/A vssd1 vssd1 vccd1 vccd1 _13738_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_32_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_231_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16457_ _16464_/B _16454_/X _16455_/X _16456_/X vssd1 vssd1 vccd1 vccd1 _18684_/D
+ sky130_fd_sc_hd__o211a_1
X_13669_ _18846_/Q _13719_/A _13752_/A _18852_/Q _13668_/X vssd1 vssd1 vccd1 vccd1
+ _13669_/X sky130_fd_sc_hd__a221o_1
XFILLER_84_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15408_ _18471_/Q _18435_/Q _15412_/S vssd1 vssd1 vccd1 vccd1 _15408_/X sky130_fd_sc_hd__mux2_1
X_19176_ _19176_/A _09008_/Y vssd1 vssd1 vccd1 vccd1 io_out[14] sky130_fd_sc_hd__ebufn_8
X_16388_ _18703_/Q _18667_/Q _16400_/S vssd1 vssd1 vccd1 vccd1 _16388_/X sky130_fd_sc_hd__mux2_1
XFILLER_191_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18127_ _19028_/CLK _18127_/D vssd1 vssd1 vccd1 vccd1 _18127_/Q sky130_fd_sc_hd__dfxtp_2
X_15339_ _15375_/A _15339_/B vssd1 vssd1 vccd1 vccd1 _15339_/Y sky130_fd_sc_hd__nand2_1
XFILLER_133_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18058_ _18069_/CLK _18058_/D vssd1 vssd1 vccd1 vccd1 _18058_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_172_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09900_ _09972_/B vssd1 vssd1 vccd1 vccd1 _10274_/S sky130_fd_sc_hd__buf_4
X_17009_ _18851_/Q _18815_/Q _17026_/S vssd1 vssd1 vccd1 vccd1 _17009_/X sky130_fd_sc_hd__mux2_1
XFILLER_67_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_1331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09831_ _11032_/A _09831_/B vssd1 vssd1 vccd1 vccd1 _12112_/C sky130_fd_sc_hd__xnor2_1
XFILLER_101_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09762_ _09764_/A _09764_/B vssd1 vssd1 vccd1 vccd1 _09816_/B sky130_fd_sc_hd__or2_1
XFILLER_6_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09693_ _10893_/S vssd1 vssd1 vccd1 vccd1 _09694_/A sky130_fd_sc_hd__buf_4
XTAP_2209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_227_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_215_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_228_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_228_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_223_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_211_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_195_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_210_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_176_wb_clk_i clkbuf_5_11_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18222_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_195_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_182_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09127_ _18842_/Q _18841_/Q _18840_/Q vssd1 vssd1 vccd1 vccd1 _09131_/A sky130_fd_sc_hd__or3_4
XFILLER_41_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_105_wb_clk_i clkbuf_5_29_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18546_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_136_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_159_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09058_ _09058_/A vssd1 vssd1 vccd1 vccd1 _09058_/Y sky130_fd_sc_hd__inv_2
XFILLER_68_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_1330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11020_ _11044_/A vssd1 vssd1 vccd1 vccd1 _13344_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_173_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_1355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_213_1352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12971_ _17985_/Q _12951_/Y _12970_/Y _12935_/X _12952_/X vssd1 vssd1 vccd1 vccd1
+ _12971_/X sky130_fd_sc_hd__o221a_1
XFILLER_66_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14710_ _14841_/B vssd1 vssd1 vccd1 vccd1 _14757_/C sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_3433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11922_ _11922_/A _11922_/B vssd1 vssd1 vccd1 vccd1 _13509_/B sky130_fd_sc_hd__xnor2_4
XFILLER_79_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_85_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15690_ _18538_/Q _18502_/Q _15693_/S vssd1 vssd1 vccd1 vccd1 _15690_/X sky130_fd_sc_hd__mux2_1
XTAP_3455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14641_ _16909_/A vssd1 vssd1 vccd1 vccd1 _15233_/B sky130_fd_sc_hd__buf_6
XTAP_3488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11853_ _11820_/A _11827_/X _11851_/X _11852_/X vssd1 vssd1 vccd1 vccd1 _11853_/X
+ sky130_fd_sc_hd__a211o_1
XTAP_2754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10804_ _09170_/A _09165_/D _09160_/D _09170_/C _10662_/A _10781_/S vssd1 vssd1 vccd1
+ vccd1 _10805_/C sky130_fd_sc_hd__mux4_2
X_17360_ _17395_/A _17360_/B vssd1 vssd1 vccd1 vccd1 _17360_/Y sky130_fd_sc_hd__nand2_1
X_14572_ _14604_/A _14574_/B vssd1 vssd1 vccd1 vccd1 _14572_/Y sky130_fd_sc_hd__nand2_1
XFILLER_25_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11784_ _11784_/A _11784_/B vssd1 vssd1 vccd1 vccd1 _11784_/X sky130_fd_sc_hd__xor2_1
XTAP_2798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_213_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16311_ _16317_/B _16309_/X _16310_/X _16295_/X vssd1 vssd1 vccd1 vccd1 _18648_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_198_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13523_ _13523_/A vssd1 vssd1 vccd1 vccd1 _13524_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_158_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10735_ _10864_/A _10833_/B _10715_/X _10725_/X _10734_/X vssd1 vssd1 vccd1 vccd1
+ _10735_/X sky130_fd_sc_hd__a311o_2
XFILLER_15_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17291_ _17336_/A _17291_/B vssd1 vssd1 vccd1 vccd1 _17291_/Y sky130_fd_sc_hd__nand2_1
XFILLER_203_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_186_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19030_ _19030_/CLK _19030_/D vssd1 vssd1 vccd1 vccd1 _19030_/Q sky130_fd_sc_hd__dfxtp_1
X_16242_ _18668_/Q _18632_/Q _16250_/S vssd1 vssd1 vccd1 vccd1 _16242_/X sky130_fd_sc_hd__mux2_1
XFILLER_186_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10666_ _10805_/A vssd1 vssd1 vccd1 vccd1 _10753_/A sky130_fd_sc_hd__buf_2
X_13454_ _13446_/Y _11655_/B _13441_/X vssd1 vssd1 vccd1 vccd1 _13455_/C sky130_fd_sc_hd__o21a_1
XFILLER_90_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12405_ _12406_/A _12406_/B _12406_/C vssd1 vssd1 vccd1 vccd1 _12414_/B sky130_fd_sc_hd__o21a_1
X_16173_ _16173_/A vssd1 vssd1 vccd1 vccd1 _16192_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_154_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13385_ _18116_/Q _11042_/X _11025_/B _11045_/X _13383_/X vssd1 vssd1 vccd1 vccd1
+ _18116_/D sky130_fd_sc_hd__o221a_1
X_10597_ _09695_/X _09696_/X _09697_/X _09698_/X _09947_/A _10307_/S vssd1 vssd1 vccd1
+ vccd1 _10598_/B sky130_fd_sc_hd__mux4_1
XFILLER_12_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15124_ _15132_/B _15121_/X _15122_/X _15123_/X vssd1 vssd1 vccd1 vccd1 _18369_/D
+ sky130_fd_sc_hd__o211a_1
X_12336_ _17889_/Q _12336_/B _12336_/C vssd1 vssd1 vccd1 vccd1 _12336_/X sky130_fd_sc_hd__or3_2
XFILLER_217_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15055_ _15061_/B _15052_/X _15054_/X _15046_/X vssd1 vssd1 vccd1 vccd1 _18351_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_141_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12267_ _12267_/A _12272_/A _12276_/C vssd1 vssd1 vccd1 vccd1 _12267_/X sky130_fd_sc_hd__and3_1
XFILLER_218_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11218_ _12940_/A vssd1 vssd1 vccd1 vccd1 _11218_/X sky130_fd_sc_hd__buf_8
X_14006_ _18946_/Q _13616_/A _13759_/A _18949_/Q _14005_/X vssd1 vssd1 vccd1 vccd1
+ _14006_/X sky130_fd_sc_hd__a221o_4
XFILLER_214_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_218_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12198_ _12198_/A _12498_/A _12198_/C vssd1 vssd1 vccd1 vccd1 _12358_/B sky130_fd_sc_hd__nor3_2
XFILLER_110_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_214_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_214_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18814_ _18823_/CLK _18814_/D vssd1 vssd1 vccd1 vccd1 _18814_/Q sky130_fd_sc_hd__dfxtp_2
X_11149_ _11764_/A _11201_/A _11149_/S vssd1 vssd1 vccd1 vccd1 _11150_/A sky130_fd_sc_hd__mux2_1
XTAP_6070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18745_ _18752_/CLK _18745_/D vssd1 vssd1 vccd1 vccd1 _18745_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_23_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15957_ _15957_/A vssd1 vssd1 vccd1 vccd1 _17228_/A sky130_fd_sc_hd__buf_8
XTAP_5391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_5_3_0_wb_clk_i clkbuf_5_3_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _17803_/CLK
+ sky130_fd_sc_hd__clkbuf_2
X_14908_ _14958_/A vssd1 vssd1 vccd1 vccd1 _14934_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_23_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18676_ _18677_/CLK _18676_/D vssd1 vssd1 vccd1 vccd1 _18676_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_149_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15888_ _18587_/Q _18551_/Q _15899_/S vssd1 vssd1 vccd1 vccd1 _15888_/X sky130_fd_sc_hd__mux2_1
XTAP_4690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17627_ _17627_/A vssd1 vssd1 vccd1 vccd1 _18969_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_224_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14839_ _14881_/A vssd1 vssd1 vccd1 vccd1 _14839_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_91_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_225_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17558_ _17548_/Y _17552_/X _18953_/Q vssd1 vssd1 vccd1 vccd1 _17558_/X sky130_fd_sc_hd__a21o_1
XFILLER_205_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_225_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_3_wb_clk_i clkbuf_5_0_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18988_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_16509_ _18734_/Q _18698_/Q _16509_/S vssd1 vssd1 vccd1 vccd1 _16509_/X sky130_fd_sc_hd__mux2_1
XFILLER_20_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_220_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17489_ _17512_/A _17489_/B vssd1 vssd1 vccd1 vccd1 _17489_/Y sky130_fd_sc_hd__nand2_1
XFILLER_220_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_225_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19228_ _19228_/A _08933_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[28] sky130_fd_sc_hd__ebufn_8
XFILLER_220_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_176_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19159_ _19159_/A _09032_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[29] sky130_fd_sc_hd__ebufn_8
XFILLER_117_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09814_ _10366_/B vssd1 vssd1 vccd1 vccd1 _12131_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_98_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_189_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09745_ _09800_/A _09800_/B vssd1 vssd1 vccd1 vccd1 _09746_/B sky130_fd_sc_hd__xor2_1
XFILLER_227_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09676_ _18239_/Q _18238_/Q _18237_/Q vssd1 vssd1 vccd1 vccd1 _09676_/X sky130_fd_sc_hd__or3_4
XTAP_2017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_210_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_1176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10520_ _10932_/A _10520_/B vssd1 vssd1 vccd1 vccd1 _10520_/X sky130_fd_sc_hd__and2_1
XFILLER_211_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_210_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_183_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10451_ _09277_/C _09277_/D _10503_/S vssd1 vssd1 vccd1 vccd1 _10451_/X sky130_fd_sc_hd__mux2_1
XFILLER_136_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13170_ _13170_/A vssd1 vssd1 vccd1 vccd1 _18042_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_201_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10382_ _10575_/A _10391_/B vssd1 vssd1 vccd1 vccd1 _10382_/X sky130_fd_sc_hd__or2_1
XFILLER_191_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12121_ _12121_/A _13526_/B vssd1 vssd1 vccd1 vccd1 _12127_/A sky130_fd_sc_hd__xnor2_1
XFILLER_151_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12052_ _12053_/A _12053_/B _13710_/A vssd1 vssd1 vccd1 vccd1 _12054_/C sky130_fd_sc_hd__a21oi_1
XFILLER_111_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11003_ _11892_/B _11237_/B _17824_/Q _11892_/A vssd1 vssd1 vccd1 vccd1 _11003_/X
+ sky130_fd_sc_hd__and4bb_1
Xclkbuf_leaf_73_wb_clk_i clkbuf_5_21_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18668_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_16860_ _16884_/A _16860_/B vssd1 vssd1 vccd1 vccd1 _16860_/Y sky130_fd_sc_hd__nand2_1
XFILLER_120_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_172_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15811_ _15857_/A _15964_/B _15811_/C vssd1 vssd1 vccd1 vccd1 _15811_/X sky130_fd_sc_hd__or3_1
X_16791_ _18803_/Q _18767_/Q _16802_/S vssd1 vssd1 vccd1 vccd1 _16791_/X sky130_fd_sc_hd__mux2_1
XFILLER_18_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_93_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18530_ _18533_/CLK _18530_/D vssd1 vssd1 vccd1 vccd1 _18530_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_20_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_218_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15742_ _18551_/Q _18515_/Q _15753_/S vssd1 vssd1 vccd1 vccd1 _15742_/X sky130_fd_sc_hd__mux2_1
XTAP_3230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12954_ _12961_/A _12949_/Y _12953_/X _12510_/X vssd1 vssd1 vccd1 vccd1 _17973_/D
+ sky130_fd_sc_hd__a211o_1
XTAP_3252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18461_ _18467_/CLK _18461_/D vssd1 vssd1 vccd1 vccd1 _18461_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_3274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11905_ _11905_/A _11973_/A vssd1 vssd1 vccd1 vccd1 _12142_/A sky130_fd_sc_hd__or2b_1
X_15673_ _15694_/A _15673_/B vssd1 vssd1 vccd1 vccd1 _15673_/Y sky130_fd_sc_hd__nand2_1
XTAP_3285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12885_ _17958_/Q _12886_/C _12884_/Y vssd1 vssd1 vccd1 vccd1 _17958_/D sky130_fd_sc_hd__a21oi_1
XTAP_2551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17412_ _17412_/A _17538_/C vssd1 vssd1 vccd1 vccd1 _17419_/B sky130_fd_sc_hd__nor2_1
X_14624_ _16886_/A vssd1 vssd1 vccd1 vccd1 _15218_/A sky130_fd_sc_hd__buf_8
XTAP_2573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18392_ _18392_/CLK _18392_/D vssd1 vssd1 vccd1 vccd1 _18392_/Q sky130_fd_sc_hd__dfxtp_2
X_11836_ _11455_/X _11470_/Y _11828_/Y vssd1 vssd1 vccd1 vccd1 _11836_/X sky130_fd_sc_hd__o21a_1
XFILLER_18_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17343_ _18934_/Q _18898_/Q _17347_/S vssd1 vssd1 vccd1 vccd1 _17343_/X sky130_fd_sc_hd__mux2_1
X_14555_ _14584_/A _14584_/B _15162_/B vssd1 vssd1 vccd1 vccd1 _14555_/X sky130_fd_sc_hd__or3_1
XTAP_1883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11767_ _11767_/A _11767_/B _11767_/C vssd1 vssd1 vccd1 vccd1 _11775_/A sky130_fd_sc_hd__and3_1
XTAP_1894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13506_ _13869_/A vssd1 vssd1 vccd1 vccd1 _13507_/A sky130_fd_sc_hd__buf_4
X_10718_ _09143_/C _09148_/B _09153_/D _09148_/D _10883_/B _10702_/A vssd1 vssd1 vccd1
+ vccd1 _10718_/X sky130_fd_sc_hd__mux4_1
X_17274_ _18880_/Q _17275_/B _17273_/Y _17260_/X vssd1 vssd1 vccd1 vccd1 _18880_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_201_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14486_ _14486_/A vssd1 vssd1 vccd1 vccd1 _18217_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_146_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11698_ _11685_/X _11709_/B _19033_/Q vssd1 vssd1 vccd1 vccd1 _11698_/X sky130_fd_sc_hd__a21bo_1
X_19013_ _19029_/CLK _19013_/D vssd1 vssd1 vccd1 vccd1 _19013_/Q sky130_fd_sc_hd__dfxtp_1
X_16225_ _16248_/A _16666_/B _16272_/C vssd1 vssd1 vccd1 vccd1 _16225_/X sky130_fd_sc_hd__or3_1
XFILLER_186_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13437_ _13438_/B _13438_/C _13438_/A vssd1 vssd1 vccd1 vccd1 _13439_/A sky130_fd_sc_hd__o21ai_1
X_10649_ _09349_/A _09354_/A _09344_/A _09349_/B _10680_/A _10648_/X vssd1 vssd1 vccd1
+ vccd1 _10649_/X sky130_fd_sc_hd__mux4_1
XFILLER_139_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16156_ _18649_/Q _18613_/Q _16170_/S vssd1 vssd1 vccd1 vccd1 _16156_/X sky130_fd_sc_hd__mux2_1
XFILLER_155_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_220_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13368_ _13368_/A _13368_/B vssd1 vssd1 vccd1 vccd1 _13368_/Y sky130_fd_sc_hd__nor2_1
XFILLER_170_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15107_ _15118_/A _15107_/B vssd1 vssd1 vccd1 vccd1 _15107_/Y sky130_fd_sc_hd__nand2_1
XFILLER_6_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12319_ _12316_/B _12329_/C _12317_/Y _12318_/X vssd1 vssd1 vccd1 vccd1 _17880_/D
+ sky130_fd_sc_hd__o211a_1
X_16087_ _18633_/Q _18597_/Q _16091_/S vssd1 vssd1 vccd1 vccd1 _16087_/X sky130_fd_sc_hd__mux2_1
XFILLER_142_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13299_ _18046_/Q _18049_/Q _18048_/Q _18051_/Q vssd1 vssd1 vccd1 vccd1 _13304_/A
+ sky130_fd_sc_hd__or4_1
XFILLER_5_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15038_ _15061_/A _15038_/B vssd1 vssd1 vccd1 vccd1 _15038_/Y sky130_fd_sc_hd__nand2_1
XFILLER_142_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_218_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_1318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_228_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_228_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16989_ _17098_/A vssd1 vssd1 vccd1 vccd1 _17078_/A sky130_fd_sc_hd__buf_2
XFILLER_68_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_209_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09530_ _09530_/A _09530_/B vssd1 vssd1 vccd1 vccd1 _09531_/B sky130_fd_sc_hd__nand2_1
X_18728_ _18732_/CLK _18728_/D vssd1 vssd1 vccd1 vccd1 _18728_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_114_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_209_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_224_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09461_ _09461_/A _18134_/D vssd1 vssd1 vccd1 vccd1 _09462_/A sky130_fd_sc_hd__or2_4
XFILLER_64_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18659_ _18662_/CLK _18659_/D vssd1 vssd1 vccd1 vccd1 _18659_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_52_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_224_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09392_ _09952_/A _09392_/B _09392_/C _09392_/D vssd1 vssd1 vccd1 vccd1 _09403_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_52_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_1340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_203_1351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_192_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19114__85 vssd1 vssd1 vccd1 vccd1 _19114__85/HI _19222_/A sky130_fd_sc_hd__conb_1
XFILLER_172_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_219_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09728_ _10895_/A _12056_/A _09728_/C _09728_/D vssd1 vssd1 vccd1 vccd1 _13410_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_228_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_227_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09659_ _13353_/A _09659_/B vssd1 vssd1 vccd1 vccd1 _12079_/A sky130_fd_sc_hd__xnor2_1
XTAP_1102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_231_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_191_wb_clk_i clkbuf_5_12_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18230_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_12670_ _17935_/Q _17932_/Q vssd1 vssd1 vccd1 vccd1 _12671_/A sky130_fd_sc_hd__xor2_1
XFILLER_151_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_231_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11621_ _11683_/A _11621_/B vssd1 vssd1 vccd1 vccd1 _11621_/Y sky130_fd_sc_hd__nand2_1
XTAP_1179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_230_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_120_wb_clk_i clkbuf_5_30_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18448_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_208_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14340_ _14533_/A vssd1 vssd1 vccd1 vccd1 _14340_/X sky130_fd_sc_hd__buf_2
X_11552_ _17867_/Q vssd1 vssd1 vccd1 vccd1 _11562_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_7_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10503_ _09119_/A _09109_/D _10503_/S vssd1 vssd1 vccd1 vccd1 _10503_/X sky130_fd_sc_hd__mux2_1
XFILLER_13_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11483_ _11508_/C _11483_/B _11483_/C vssd1 vssd1 vccd1 vccd1 _11484_/B sky130_fd_sc_hd__and3_1
X_14271_ _14202_/X _14268_/X _14269_/X _14270_/X vssd1 vssd1 vccd1 vccd1 _18173_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_195_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16010_ _18616_/Q _18580_/Q _16010_/S vssd1 vssd1 vccd1 vccd1 _16010_/X sky130_fd_sc_hd__mux2_1
XFILLER_143_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10434_ _10431_/X _10432_/X _10926_/A vssd1 vssd1 vccd1 vccd1 _10434_/X sky130_fd_sc_hd__mux2_2
X_13222_ _13222_/A _18067_/Q vssd1 vssd1 vccd1 vccd1 _13223_/A sky130_fd_sc_hd__and2_1
XFILLER_10_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_1266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10365_ _09889_/A _10361_/X _10364_/X _12126_/A vssd1 vssd1 vccd1 vccd1 _10365_/X
+ sky130_fd_sc_hd__a22o_1
X_13153_ _13153_/A input3/X vssd1 vssd1 vccd1 vccd1 _18035_/D sky130_fd_sc_hd__nor2_1
XFILLER_152_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12104_ _12104_/A _12104_/B _12104_/C _12104_/D vssd1 vssd1 vccd1 vccd1 _12104_/X
+ sky130_fd_sc_hd__or4_1
XFILLER_112_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13084_ _17420_/A vssd1 vssd1 vccd1 vccd1 _14480_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_17961_ _17965_/CLK _17961_/D vssd1 vssd1 vccd1 vccd1 _17961_/Q sky130_fd_sc_hd__dfxtp_1
X_10296_ _10291_/X _10292_/X _10295_/X _10370_/S vssd1 vssd1 vccd1 vccd1 _10296_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_124_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_215_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16912_ _18829_/Q _18793_/Q _16925_/S vssd1 vssd1 vccd1 vccd1 _16912_/X sky130_fd_sc_hd__mux2_1
X_12035_ _11924_/Y _11925_/X _11993_/X _12034_/X vssd1 vssd1 vccd1 vccd1 _12035_/X
+ sky130_fd_sc_hd__a211o_1
X_17892_ _17895_/CLK _17892_/D vssd1 vssd1 vccd1 vccd1 _17892_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_214_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16843_ _16882_/A _16847_/B vssd1 vssd1 vccd1 vccd1 _16843_/Y sky130_fd_sc_hd__nand2_1
XFILLER_78_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_219_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16774_ _16779_/B _16772_/X _16773_/X _16760_/X vssd1 vssd1 vccd1 vccd1 _18762_/D
+ sky130_fd_sc_hd__o211a_1
X_13986_ _18406_/Q _13613_/A _13670_/X _18400_/Q vssd1 vssd1 vccd1 vccd1 _13986_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_20_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_1351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18513_ _18548_/CLK _18513_/D vssd1 vssd1 vccd1 vccd1 _18513_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_59_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_1362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15725_ _15730_/B _15723_/X _15724_/X _15720_/X vssd1 vssd1 vccd1 vccd1 _18510_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_18_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12937_ _11031_/A _11036_/B _12935_/X _12933_/A _12936_/Y vssd1 vssd1 vccd1 vccd1
+ _12939_/A sky130_fd_sc_hd__o311a_1
XFILLER_185_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_208_wb_clk_i _17803_/CLK vssd1 vssd1 vccd1 vccd1 _18972_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_3071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_207_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_222_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18444_ _18448_/CLK _18444_/D vssd1 vssd1 vccd1 vccd1 _18444_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_33_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15656_ _15661_/B _15654_/X _15655_/X _15640_/X vssd1 vssd1 vccd1 vccd1 _18492_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_179_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_1338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12868_ _17953_/Q _12868_/B vssd1 vssd1 vccd1 vccd1 _12869_/A sky130_fd_sc_hd__and2_1
XFILLER_15_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_222_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14607_ _18245_/Q _14606_/B _14606_/Y _14587_/X vssd1 vssd1 vccd1 vccd1 _18245_/D
+ sky130_fd_sc_hd__o211a_1
X_18375_ _18380_/CLK _18375_/D vssd1 vssd1 vccd1 vccd1 _18375_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_33_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11819_ _11742_/X _11778_/X _11818_/Y _11809_/X vssd1 vssd1 vccd1 vccd1 _11820_/B
+ sky130_fd_sc_hd__a31o_1
X_15587_ _15613_/A _16032_/B _15599_/C vssd1 vssd1 vccd1 vccd1 _15587_/X sky130_fd_sc_hd__or3_1
XFILLER_33_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12799_ _17954_/Q vssd1 vssd1 vccd1 vccd1 _12871_/A sky130_fd_sc_hd__inv_2
XFILLER_14_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17326_ _18929_/Q _18893_/Q _17347_/S vssd1 vssd1 vccd1 vccd1 _17326_/X sky130_fd_sc_hd__mux2_1
X_14538_ _17541_/A vssd1 vssd1 vccd1 vccd1 _14604_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_175_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_222_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17257_ _17263_/B _17255_/X _17256_/X _17241_/X vssd1 vssd1 vccd1 vccd1 _18876_/D
+ sky130_fd_sc_hd__o211a_1
X_14469_ _14470_/B _14464_/A _14464_/B _14470_/A vssd1 vssd1 vccd1 vccd1 _14471_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_128_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16208_ _16248_/A _16796_/B _16208_/C vssd1 vssd1 vccd1 vccd1 _16208_/X sky130_fd_sc_hd__or3_1
XFILLER_134_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17188_ _18859_/Q _17189_/B _17187_/Y _17181_/X vssd1 vssd1 vccd1 vccd1 _18859_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_115_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16139_ _16139_/A vssd1 vssd1 vccd1 vccd1 _16139_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_192_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_170_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08961_ _08967_/A vssd1 vssd1 vccd1 vccd1 _08966_/A sky130_fd_sc_hd__buf_12
XFILLER_192_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_190_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_217_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09513_ _18230_/Q _18229_/Q _18228_/Q vssd1 vssd1 vccd1 vccd1 _14372_/B sky130_fd_sc_hd__or3_1
XFILLER_83_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_225_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_213_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_225_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_213_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09444_ _09450_/B _09441_/X _09442_/X _09443_/Y vssd1 vssd1 vccd1 vccd1 _09444_/Y
+ sky130_fd_sc_hd__o211ai_4
XFILLER_25_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_224_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_220_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_212_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09375_ _18386_/Q _18385_/Q _18384_/Q vssd1 vssd1 vccd1 vccd1 _09376_/D sky130_fd_sc_hd__or3_4
XFILLER_36_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_192_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_181_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10150_ _19027_/Q vssd1 vssd1 vccd1 vccd1 _10155_/A sky130_fd_sc_hd__clkbuf_2
XTAP_5902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10081_ _09657_/A _10077_/X _10080_/X _09720_/X vssd1 vssd1 vccd1 vccd1 _10081_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_5924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_181_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13840_ _18682_/Q _13524_/A _14026_/A _18688_/Q vssd1 vssd1 vccd1 vccd1 _13840_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_74_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_216_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_210_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13771_ _12027_/C _13757_/X _13770_/X _12028_/A vssd1 vssd1 vccd1 vccd1 _13829_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_43_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10983_ _18996_/Q vssd1 vssd1 vccd1 vccd1 _14187_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_15510_ _18494_/Q _18458_/Q _15514_/S vssd1 vssd1 vccd1 vccd1 _15510_/X sky130_fd_sc_hd__mux2_1
XFILLER_43_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12722_ _18088_/Q vssd1 vssd1 vccd1 vccd1 _12925_/B sky130_fd_sc_hd__inv_2
X_16490_ _18729_/Q _18693_/Q _16490_/S vssd1 vssd1 vccd1 vccd1 _16490_/X sky130_fd_sc_hd__mux2_1
XFILLER_31_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15441_ _18478_/Q _18442_/Q _15458_/S vssd1 vssd1 vccd1 vccd1 _15441_/X sky130_fd_sc_hd__mux2_1
XFILLER_130_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12653_ _17933_/Q _12653_/B vssd1 vssd1 vccd1 vccd1 _12654_/B sky130_fd_sc_hd__and2_1
XFILLER_145_1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11604_ _17857_/Q vssd1 vssd1 vccd1 vccd1 _12233_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_30_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18160_ _18163_/CLK _18160_/D vssd1 vssd1 vccd1 vccd1 _18160_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_54_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15372_ _18426_/Q _15375_/B _15371_/X _15363_/X vssd1 vssd1 vccd1 vccd1 _18426_/D
+ sky130_fd_sc_hd__o211a_1
X_12584_ _12582_/A _12582_/B _12613_/A vssd1 vssd1 vccd1 vccd1 _12584_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_180_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17111_ _18877_/Q _18841_/Q _17114_/S vssd1 vssd1 vccd1 vccd1 _17111_/X sky130_fd_sc_hd__mux2_1
X_14323_ _18208_/Q _14323_/B _14323_/C vssd1 vssd1 vccd1 vccd1 _14325_/A sky130_fd_sc_hd__or3_1
XFILLER_156_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11535_ _12279_/A _11390_/A _11531_/Y _11534_/Y _11619_/A vssd1 vssd1 vccd1 vccd1
+ _11535_/X sky130_fd_sc_hd__o32a_1
X_18091_ _18224_/CLK _18091_/D vssd1 vssd1 vccd1 vccd1 _18091_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_184_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_221_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17042_ _17164_/A vssd1 vssd1 vccd1 vccd1 _17088_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_116_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14254_ _14243_/X _14227_/X _14229_/X _14244_/X _18171_/Q vssd1 vssd1 vccd1 vccd1
+ _14254_/X sky130_fd_sc_hd__a311o_1
XFILLER_137_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11466_ _11586_/A _11466_/B vssd1 vssd1 vccd1 vccd1 _11593_/A sky130_fd_sc_hd__nand2_2
XFILLER_109_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13205_ _13205_/A vssd1 vssd1 vccd1 vccd1 _18058_/D sky130_fd_sc_hd__clkbuf_1
X_10417_ _10932_/A vssd1 vssd1 vccd1 vccd1 _10419_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_11397_ _11541_/A _11541_/B vssd1 vssd1 vccd1 vccd1 _11542_/B sky130_fd_sc_hd__or2_1
X_14185_ _14185_/A _14185_/B vssd1 vssd1 vccd1 vccd1 _18168_/D sky130_fd_sc_hd__nand2_1
XFILLER_174_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_124_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13136_ _13140_/A _18028_/Q vssd1 vssd1 vccd1 vccd1 _13137_/A sky130_fd_sc_hd__and2_1
XTAP_705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10348_ _10348_/A vssd1 vssd1 vccd1 vccd1 _10349_/S sky130_fd_sc_hd__buf_6
XFILLER_225_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18993_ _18993_/CLK _18993_/D vssd1 vssd1 vccd1 vccd1 _18993_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10279_ _09181_/B _09176_/C _10286_/S vssd1 vssd1 vccd1 vccd1 _10279_/X sky130_fd_sc_hd__mux2_1
XTAP_749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17944_ _18213_/CLK _17944_/D vssd1 vssd1 vccd1 vccd1 _17944_/Q sky130_fd_sc_hd__dfxtp_2
X_13067_ _13067_/A vssd1 vssd1 vccd1 vccd1 _17999_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_215_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12018_ _12018_/A _12049_/B vssd1 vssd1 vccd1 vccd1 _12019_/B sky130_fd_sc_hd__nor2_8
XFILLER_22_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17875_ _17879_/CLK _17875_/D vssd1 vssd1 vccd1 vccd1 _17875_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_78_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_113_1326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_227_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16826_ _16833_/B _16822_/X _16824_/X _16825_/X vssd1 vssd1 vccd1 vccd1 _18774_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_65_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16757_ _16757_/A _16794_/B vssd1 vssd1 vccd1 vccd1 _16769_/B sky130_fd_sc_hd__nor2_2
X_13969_ _18445_/Q _13759_/X _13780_/X _18436_/Q _13968_/X vssd1 vssd1 vccd1 vccd1
+ _13969_/X sky130_fd_sc_hd__a221o_4
XFILLER_19_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15708_ _15754_/A _15708_/B vssd1 vssd1 vccd1 vccd1 _15708_/Y sky130_fd_sc_hd__nand2_1
XFILLER_146_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16688_ _16727_/A vssd1 vssd1 vccd1 vccd1 _16745_/B sky130_fd_sc_hd__buf_2
XFILLER_55_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_206_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18427_ _18434_/CLK _18427_/D vssd1 vssd1 vccd1 vccd1 _18427_/Q sky130_fd_sc_hd__dfxtp_1
X_15639_ _15739_/A vssd1 vssd1 vccd1 vccd1 _15720_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_146_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_107_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09160_ _09160_/A _09160_/B _09160_/C _09160_/D vssd1 vssd1 vccd1 vccd1 _09171_/A
+ sky130_fd_sc_hd__and4_1
X_18358_ _18387_/CLK _18358_/D vssd1 vssd1 vccd1 vccd1 _18358_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_222_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_202_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17309_ _17314_/B _17307_/X _17308_/X _17304_/X vssd1 vssd1 vccd1 vccd1 _18888_/D
+ sky130_fd_sc_hd__o211a_1
X_09091_ _18776_/Q _18775_/Q _18774_/Q vssd1 vssd1 vccd1 vccd1 _09093_/C sky130_fd_sc_hd__or3_4
XFILLER_119_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18289_ _18290_/CLK _18289_/D vssd1 vssd1 vccd1 vccd1 _18289_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_190_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09993_ _09993_/A _10004_/B vssd1 vssd1 vccd1 vccd1 _09993_/X sky130_fd_sc_hd__or2_1
XFILLER_135_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08944_ _08948_/A vssd1 vssd1 vccd1 vccd1 _08944_/Y sky130_fd_sc_hd__inv_2
XFILLER_131_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_151_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_217_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_217_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_226_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_212_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09427_ _09427_/A _09427_/B vssd1 vssd1 vccd1 vccd1 _09427_/Y sky130_fd_sc_hd__nand2_1
XFILLER_52_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_213_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_197_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_212_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_139_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09358_ _18275_/Q _18274_/Q _18273_/Q vssd1 vssd1 vccd1 vccd1 _09360_/C sky130_fd_sc_hd__or3_2
XFILLER_100_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09289_ _09435_/A _09432_/C vssd1 vssd1 vccd1 vccd1 _09454_/B sky130_fd_sc_hd__and2b_1
XFILLER_193_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11320_ _17876_/Q vssd1 vssd1 vccd1 vccd1 _11345_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_138_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11251_ _11405_/A vssd1 vssd1 vccd1 vccd1 _11735_/B sky130_fd_sc_hd__buf_2
XFILLER_10_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_180_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10202_ _10202_/A _10202_/B vssd1 vssd1 vccd1 vccd1 _10217_/B sky130_fd_sc_hd__or2_1
XFILLER_136_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11182_ _11185_/B _11198_/B _11182_/C vssd1 vssd1 vccd1 vccd1 _11183_/A sky130_fd_sc_hd__and3b_1
XFILLER_69_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_1348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10133_ _10133_/A vssd1 vssd1 vccd1 vccd1 _10146_/A sky130_fd_sc_hd__inv_2
XFILLER_69_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15990_ _18611_/Q _18575_/Q _15990_/S vssd1 vssd1 vccd1 vccd1 _15990_/X sky130_fd_sc_hd__mux2_1
XTAP_5721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14941_ _14980_/A vssd1 vssd1 vccd1 vccd1 _14941_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_10064_ _09176_/C _10008_/A _10063_/X vssd1 vssd1 vccd1 vccd1 _10065_/C sky130_fd_sc_hd__a21o_1
XTAP_5754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17660_ _17660_/A vssd1 vssd1 vccd1 vccd1 _18977_/D sky130_fd_sc_hd__clkbuf_1
XTAP_5798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14872_ _14872_/A _14875_/B vssd1 vssd1 vccd1 vccd1 _14872_/Y sky130_fd_sc_hd__nand2_1
XFILLER_63_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16611_ _16634_/A _16611_/B vssd1 vssd1 vccd1 vccd1 _16611_/Y sky130_fd_sc_hd__nand2_1
XFILLER_76_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13823_ _18573_/Q _13785_/A _13535_/A _18555_/Q vssd1 vssd1 vccd1 vccd1 _13823_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_90_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17591_ _17591_/A vssd1 vssd1 vccd1 vccd1 _17591_/X sky130_fd_sc_hd__clkbuf_2
XINSDIODE2_106 _13940_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINSDIODE2_117 _16839_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16542_ _16689_/A _16602_/B vssd1 vssd1 vccd1 vccd1 _16551_/B sky130_fd_sc_hd__nor2_1
XINSDIODE2_128 _16219_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13754_ _18795_/Q _13529_/A _13725_/X _18771_/Q vssd1 vssd1 vccd1 vccd1 _13754_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_56_1305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XINSDIODE2_139 _15440_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10966_ _12056_/A _10966_/B vssd1 vssd1 vccd1 vccd1 _10966_/Y sky130_fd_sc_hd__nand2_1
XFILLER_16_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12705_ _17936_/Q _12523_/X _12704_/X _12510_/X vssd1 vssd1 vccd1 vccd1 _17936_/D
+ sky130_fd_sc_hd__a211o_1
X_16473_ _16473_/A vssd1 vssd1 vccd1 vccd1 _16490_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_204_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13685_ _13731_/A vssd1 vssd1 vccd1 vccd1 _13697_/A sky130_fd_sc_hd__buf_4
X_10897_ _10897_/A _10897_/B _10897_/C _10896_/Y vssd1 vssd1 vccd1 vccd1 _10897_/X
+ sky130_fd_sc_hd__or4b_1
X_18212_ _18213_/CLK _18212_/D vssd1 vssd1 vccd1 vccd1 _18212_/Q sky130_fd_sc_hd__dfxtp_1
X_15424_ _15431_/B _15421_/X _15423_/X _15404_/X vssd1 vssd1 vccd1 vccd1 _18438_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_148_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_188_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19192_ _19192_/A _08993_/Y vssd1 vssd1 vccd1 vccd1 io_out[30] sky130_fd_sc_hd__ebufn_8
X_12636_ _17931_/Q _12637_/B vssd1 vssd1 vccd1 vccd1 _12638_/A sky130_fd_sc_hd__nor2_1
XFILLER_223_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18143_ _18147_/CLK _18143_/D vssd1 vssd1 vccd1 vccd1 _18143_/Q sky130_fd_sc_hd__dfxtp_1
X_15355_ _15962_/A _15393_/B vssd1 vssd1 vccd1 vccd1 _15366_/B sky130_fd_sc_hd__nor2_2
XFILLER_200_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12567_ _12561_/Y _12563_/Y _12565_/X _12635_/A vssd1 vssd1 vccd1 vccd1 _12567_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_145_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14306_ _14464_/A _14305_/A _14335_/B _14305_/Y vssd1 vssd1 vccd1 vccd1 _14306_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_184_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11518_ _17872_/Q _17871_/Q _17870_/Q vssd1 vssd1 vccd1 vccd1 _12287_/A sky130_fd_sc_hd__nand3_1
X_18074_ _18085_/CLK _18074_/D vssd1 vssd1 vccd1 vccd1 _18074_/Q sky130_fd_sc_hd__dfxtp_1
X_15286_ _15303_/A _15286_/B vssd1 vssd1 vccd1 vccd1 _15286_/Y sky130_fd_sc_hd__nand2_1
XFILLER_102_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12498_ _12498_/A vssd1 vssd1 vccd1 vccd1 _12498_/Y sky130_fd_sc_hd__inv_2
XFILLER_171_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17025_ _17458_/A _17070_/B vssd1 vssd1 vccd1 vccd1 _17035_/B sky130_fd_sc_hd__nor2_2
XFILLER_116_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14237_ _14237_/A vssd1 vssd1 vccd1 vccd1 _14237_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_144_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11449_ _13485_/A _11442_/A _11654_/C _11922_/A vssd1 vssd1 vccd1 vccd1 _11496_/A
+ sky130_fd_sc_hd__a31o_1
XFILLER_171_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14168_ _18608_/Q _13568_/A _13515_/A _18602_/Q vssd1 vssd1 vccd1 vccd1 _14168_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_124_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13119_ _13119_/A vssd1 vssd1 vccd1 vccd1 _18019_/D sky130_fd_sc_hd__clkbuf_1
XTAP_524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14099_ _18632_/Q _14019_/A _13500_/A _18656_/Q vssd1 vssd1 vccd1 vccd1 _14099_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18976_ _18977_/CLK _18976_/D vssd1 vssd1 vccd1 vccd1 _18976_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_230_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17927_ _17931_/CLK _17927_/D vssd1 vssd1 vccd1 vccd1 _17927_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_223_wb_clk_i _17803_/CLK vssd1 vssd1 vccd1 vccd1 _18191_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_227_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_230_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_227_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17858_ _17861_/CLK _17858_/D vssd1 vssd1 vccd1 vccd1 _17858_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_82_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16809_ _16879_/A vssd1 vssd1 vccd1 vccd1 _16960_/B sky130_fd_sc_hd__buf_2
XFILLER_81_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17789_ _17793_/CLK _17789_/D vssd1 vssd1 vccd1 vccd1 _17789_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_198_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_223_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_224_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_222_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_222_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09212_ _18668_/Q _18667_/Q _18666_/Q vssd1 vssd1 vccd1 vccd1 _09214_/C sky130_fd_sc_hd__or3_4
XFILLER_22_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09143_ _09993_/A _09143_/B _09143_/C _09143_/D vssd1 vssd1 vccd1 vccd1 _09154_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_147_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09074_ _17838_/Q vssd1 vssd1 vccd1 vccd1 _09083_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_163_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09976_ _09976_/A vssd1 vssd1 vccd1 vccd1 _10605_/B sky130_fd_sc_hd__buf_4
XTAP_5017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_229_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10820_ _13007_/A _10820_/B vssd1 vssd1 vccd1 vccd1 _10821_/B sky130_fd_sc_hd__nor2_2
XTAP_2947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_213_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_98_wb_clk_i clkbuf_5_28_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18149_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_10751_ _10679_/X _10735_/X _10750_/X _10678_/X vssd1 vssd1 vccd1 vccd1 _10752_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_198_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13470_ _17843_/Q _13457_/X _13465_/X vssd1 vssd1 vccd1 vccd1 _13471_/B sky130_fd_sc_hd__a21oi_1
Xclkbuf_leaf_27_wb_clk_i clkbuf_5_7_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18939_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_231_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10682_ _10701_/A vssd1 vssd1 vccd1 vccd1 _10809_/A sky130_fd_sc_hd__buf_2
XFILLER_201_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12421_ _12439_/A _12420_/X _12412_/A _12413_/X vssd1 vssd1 vccd1 vccd1 _12423_/B
+ sky130_fd_sc_hd__a211o_1
XFILLER_138_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_1268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15140_ _15142_/B _15138_/X _15139_/Y _15123_/X vssd1 vssd1 vccd1 vccd1 _18373_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_138_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12352_ _17892_/Q _12352_/B _12499_/C vssd1 vssd1 vccd1 vccd1 _12353_/A sky130_fd_sc_hd__or3_1
XFILLER_138_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11303_ _11303_/A _11635_/A _11770_/A vssd1 vssd1 vccd1 vccd1 _11842_/A sky130_fd_sc_hd__nor3b_2
XFILLER_14_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15071_ _15252_/A vssd1 vssd1 vccd1 vccd1 _15118_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_4_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12283_ _17873_/Q _12279_/A _12279_/B vssd1 vssd1 vccd1 vccd1 _12304_/B sky130_fd_sc_hd__a21oi_2
X_14022_ _18869_/Q _13532_/A _13539_/A _18845_/Q vssd1 vssd1 vccd1 vccd1 _14022_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_107_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_181_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11234_ _11234_/A _11234_/B vssd1 vssd1 vccd1 vccd1 _17820_/D sky130_fd_sc_hd__nor2_1
XFILLER_101_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_106_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_214_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_175_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18830_ _18849_/CLK _18830_/D vssd1 vssd1 vccd1 vccd1 _18830_/Q sky130_fd_sc_hd__dfxtp_2
X_11165_ _17805_/Q _11212_/B vssd1 vssd1 vccd1 vccd1 _11177_/B sky130_fd_sc_hd__and2_1
XFILLER_96_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19075__46 vssd1 vssd1 vccd1 vccd1 _19075__46/HI _19169_/A sky130_fd_sc_hd__conb_1
XFILLER_1_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10116_ _18119_/Q _10116_/B vssd1 vssd1 vccd1 vccd1 _10142_/B sky130_fd_sc_hd__xnor2_1
X_15973_ _15971_/B _15970_/X _15971_/Y _15972_/X vssd1 vssd1 vccd1 vccd1 _18569_/D
+ sky130_fd_sc_hd__o211a_1
X_18761_ _18764_/CLK _18761_/D vssd1 vssd1 vccd1 vccd1 _18761_/Q sky130_fd_sc_hd__dfxtp_2
X_11096_ _11096_/A vssd1 vssd1 vccd1 vccd1 _17793_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_62_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_212_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14924_ _14935_/A _14924_/B vssd1 vssd1 vccd1 vccd1 _14924_/Y sky130_fd_sc_hd__nand2_1
X_10047_ _09214_/A _09219_/C _09219_/D _09209_/B _10004_/B _10090_/S vssd1 vssd1 vccd1
+ vccd1 _10047_/X sky130_fd_sc_hd__mux4_1
XFILLER_23_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17712_ _17712_/A _19002_/Q vssd1 vssd1 vccd1 vccd1 _17713_/A sky130_fd_sc_hd__and2_1
XFILLER_76_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_212_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_222_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18692_ _18693_/CLK _18692_/D vssd1 vssd1 vccd1 vccd1 _18692_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_4850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14855_ _14985_/B vssd1 vssd1 vccd1 vccd1 _14906_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_17643_ _17659_/A _17643_/B vssd1 vssd1 vccd1 vccd1 _17644_/A sky130_fd_sc_hd__and2_1
XTAP_4894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_223_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13806_ _18396_/Q _13716_/X _13654_/A _18387_/Q _13805_/X vssd1 vssd1 vccd1 vccd1
+ _13806_/X sky130_fd_sc_hd__a221o_1
X_17574_ _17574_/A vssd1 vssd1 vccd1 vccd1 _18956_/D sky130_fd_sc_hd__clkbuf_1
X_14786_ _14788_/B _14784_/X _14785_/Y _14778_/X vssd1 vssd1 vccd1 vccd1 _18286_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_223_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11998_ _12041_/C _11929_/X _11997_/Y _12015_/A vssd1 vssd1 vccd1 vccd1 _12006_/A
+ sky130_fd_sc_hd__o31a_1
XFILLER_90_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16525_ _16575_/A _16525_/B vssd1 vssd1 vccd1 vccd1 _16525_/Y sky130_fd_sc_hd__nand2_1
XFILLER_56_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_220_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13737_ _18312_/Q _13734_/X _13592_/A _18330_/Q _13736_/X vssd1 vssd1 vccd1 vccd1
+ _13737_/X sky130_fd_sc_hd__a221o_1
XFILLER_108_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10949_ _10946_/X _10947_/X _10948_/X _10010_/X _09689_/X vssd1 vssd1 vccd1 vccd1
+ _10949_/X sky130_fd_sc_hd__a221o_1
XFILLER_44_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_176_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16456_ _16456_/A vssd1 vssd1 vccd1 vccd1 _16456_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_56_1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13668_ _18855_/Q _13652_/A _13720_/A _18870_/Q vssd1 vssd1 vccd1 vccd1 _13668_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_231_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15407_ _16005_/A _15448_/B vssd1 vssd1 vccd1 vccd1 _15417_/B sky130_fd_sc_hd__nor2_2
XPHY_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19175_ _19175_/A _09007_/Y vssd1 vssd1 vccd1 vccd1 io_out[13] sky130_fd_sc_hd__ebufn_8
X_12619_ _12619_/A _12619_/B vssd1 vssd1 vccd1 vccd1 _12619_/X sky130_fd_sc_hd__or2_1
X_16387_ _16392_/B _16384_/X _16386_/X _16376_/X vssd1 vssd1 vccd1 vccd1 _18666_/D
+ sky130_fd_sc_hd__o211a_1
X_13599_ _18717_/Q _13596_/X _13598_/X _18699_/Q vssd1 vssd1 vccd1 vccd1 _13599_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_118_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18126_ _18126_/CLK _18126_/D vssd1 vssd1 vccd1 vccd1 _18126_/Q sky130_fd_sc_hd__dfxtp_4
X_15338_ _18455_/Q _18419_/Q _15356_/S vssd1 vssd1 vccd1 vccd1 _15338_/X sky130_fd_sc_hd__mux2_1
X_18057_ _18069_/CLK _18057_/D vssd1 vssd1 vccd1 vccd1 _18057_/Q sky130_fd_sc_hd__dfxtp_1
X_15269_ _15275_/B _15267_/X _15268_/X _15264_/X vssd1 vssd1 vccd1 vccd1 _18405_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_144_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17008_ _17078_/A vssd1 vssd1 vccd1 vccd1 _17026_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_104_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_1264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09830_ _17976_/Q _17781_/Q vssd1 vssd1 vccd1 vccd1 _09831_/B sky130_fd_sc_hd__xnor2_1
XFILLER_112_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_1207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09761_ _09784_/A _09784_/B _09760_/X vssd1 vssd1 vccd1 vccd1 _09764_/B sky130_fd_sc_hd__o21a_1
XFILLER_39_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18959_ _18959_/CLK _18959_/D vssd1 vssd1 vccd1 vccd1 _18959_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_189_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_227_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09692_ _09692_/A _09719_/B vssd1 vssd1 vccd1 vccd1 _10893_/S sky130_fd_sc_hd__xnor2_4
XFILLER_132_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_228_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09126_ _09126_/A _09126_/B _09126_/C _09126_/D vssd1 vssd1 vccd1 vccd1 _09137_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_148_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_159_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_191_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09057_ _09058_/A vssd1 vssd1 vccd1 vccd1 _09057_/Y sky130_fd_sc_hd__inv_2
XFILLER_159_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_145_wb_clk_i clkbuf_5_26_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18296_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_2_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_1334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_1367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_106_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09959_ _09959_/A vssd1 vssd1 vccd1 vccd1 _09959_/X sky130_fd_sc_hd__buf_4
XTAP_4102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_218_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12970_ _12970_/A _12970_/B vssd1 vssd1 vccd1 vccd1 _12970_/Y sky130_fd_sc_hd__nor2_1
XFILLER_218_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11921_ _13501_/A _11921_/B vssd1 vssd1 vccd1 vccd1 _11922_/B sky130_fd_sc_hd__and2_2
XTAP_4179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14640_ _16905_/A vssd1 vssd1 vccd1 vccd1 _16909_/A sky130_fd_sc_hd__buf_4
XTAP_3478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11852_ _11867_/A vssd1 vssd1 vccd1 vccd1 _11852_/X sky130_fd_sc_hd__clkbuf_2
XTAP_2744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10803_ _09214_/A _09219_/C _09219_/D _09209_/B _10877_/B _10809_/A vssd1 vssd1 vccd1
+ vccd1 _10803_/X sky130_fd_sc_hd__mux4_2
XTAP_2777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14571_ _18237_/Q _14574_/B _14570_/X _14561_/X vssd1 vssd1 vccd1 vccd1 _18237_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_14_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11783_ _11783_/A _11783_/B vssd1 vssd1 vccd1 vccd1 _11783_/Y sky130_fd_sc_hd__nor2_1
XTAP_2799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16310_ _16310_/A _16749_/B _16333_/C vssd1 vssd1 vccd1 vccd1 _16310_/X sky130_fd_sc_hd__or3_1
XFILLER_41_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13522_ _13522_/A vssd1 vssd1 vccd1 vccd1 _13523_/A sky130_fd_sc_hd__buf_4
XFILLER_198_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_159_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10734_ _10753_/A _10726_/X _10730_/X _10733_/X vssd1 vssd1 vccd1 vccd1 _10734_/X
+ sky130_fd_sc_hd__o211a_1
X_17290_ _17468_/A vssd1 vssd1 vccd1 vccd1 _17336_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_158_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_201_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16241_ _16243_/B _16239_/X _16240_/Y _16230_/X vssd1 vssd1 vccd1 vccd1 _18631_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_186_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13453_ _13446_/Y _11655_/B _13441_/X _13451_/X _13452_/Y vssd1 vssd1 vccd1 vccd1
+ _13455_/B sky130_fd_sc_hd__o311a_1
XFILLER_55_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10665_ _09344_/C _09344_/D _09354_/D _09349_/D _10660_/X _10859_/S vssd1 vssd1 vccd1
+ vccd1 _10665_/X sky130_fd_sc_hd__mux4_2
XFILLER_167_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12404_ _12414_/A _12404_/B vssd1 vssd1 vccd1 vccd1 _12406_/C sky130_fd_sc_hd__nor2_1
X_16172_ _16175_/B _16170_/X _16171_/Y _16162_/X vssd1 vssd1 vccd1 vccd1 _18616_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_142_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_220_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13384_ _18115_/Q _11042_/X _11044_/B _11026_/A _13383_/X vssd1 vssd1 vccd1 vccd1
+ _18115_/D sky130_fd_sc_hd__o221a_1
X_10596_ _10579_/X _10585_/X _10594_/X _10110_/Y _10595_/X vssd1 vssd1 vccd1 vccd1
+ _10897_/B sky130_fd_sc_hd__o311a_1
X_15123_ _15187_/A vssd1 vssd1 vccd1 vccd1 _15123_/X sky130_fd_sc_hd__clkbuf_2
X_12335_ _17884_/Q _11431_/B _12317_/Y vssd1 vssd1 vccd1 vccd1 _12336_/C sky130_fd_sc_hd__o21bai_1
XFILLER_86_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15054_ _15098_/A _15199_/B _15054_/C vssd1 vssd1 vccd1 vccd1 _15054_/X sky130_fd_sc_hd__or3_1
XFILLER_147_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12266_ _12269_/B _12269_/C _12270_/B vssd1 vssd1 vccd1 vccd1 _12266_/X sky130_fd_sc_hd__and3_1
XFILLER_107_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_218_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14005_ _18922_/Q _13733_/A _14001_/X _14004_/X vssd1 vssd1 vccd1 vccd1 _14005_/X
+ sky130_fd_sc_hd__a211o_1
X_11217_ _16891_/A vssd1 vssd1 vccd1 vccd1 _12940_/A sky130_fd_sc_hd__clkbuf_2
X_12197_ _17900_/Q _17899_/Q _12197_/C _12476_/B vssd1 vssd1 vccd1 vccd1 _12198_/C
+ sky130_fd_sc_hd__or4_1
XFILLER_218_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18813_ _18823_/CLK _18813_/D vssd1 vssd1 vccd1 vccd1 _18813_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_122_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_96_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11148_ _11770_/A vssd1 vssd1 vccd1 vccd1 _11764_/A sky130_fd_sc_hd__buf_2
XTAP_6071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_209_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18744_ _18752_/CLK _18744_/D vssd1 vssd1 vccd1 vccd1 _18744_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_62_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15956_ _18602_/Q _18566_/Q _15963_/S vssd1 vssd1 vccd1 vccd1 _15956_/X sky130_fd_sc_hd__mux2_1
XTAP_5370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11079_ _17790_/Q vssd1 vssd1 vccd1 vccd1 _11970_/A sky130_fd_sc_hd__clkbuf_2
XTAP_5381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14907_ _14913_/B _14905_/X _14906_/X _14902_/X vssd1 vssd1 vccd1 vccd1 _18315_/D
+ sky130_fd_sc_hd__o211a_1
X_18675_ _18677_/CLK _18675_/D vssd1 vssd1 vccd1 vccd1 _18675_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_209_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15887_ _15890_/B _15884_/X _15886_/Y _15881_/X vssd1 vssd1 vccd1 vccd1 _18550_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_4680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17626_ _17638_/A _17626_/B vssd1 vssd1 vccd1 vccd1 _17627_/A sky130_fd_sc_hd__and2_1
X_14838_ _14875_/A _14838_/B vssd1 vssd1 vccd1 vccd1 _14838_/Y sky130_fd_sc_hd__nand2_1
XFILLER_149_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_225_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17557_ _14357_/X _16975_/X _17547_/X _17555_/X _17556_/X vssd1 vssd1 vccd1 vccd1
+ _18952_/D sky130_fd_sc_hd__o311a_1
X_14769_ _14915_/A vssd1 vssd1 vccd1 vccd1 _17473_/B sky130_fd_sc_hd__buf_8
XFILLER_205_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16508_ _16510_/B _16506_/X _16507_/Y _16496_/X vssd1 vssd1 vccd1 vccd1 _18697_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_225_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17488_ _18971_/Q _18935_/Q _17495_/S vssd1 vssd1 vccd1 vccd1 _17488_/X sky130_fd_sc_hd__mux2_1
XFILLER_149_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19227_ _19227_/A _08934_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[27] sky130_fd_sc_hd__ebufn_8
X_16439_ _16450_/A _16439_/B vssd1 vssd1 vccd1 vccd1 _16439_/Y sky130_fd_sc_hd__nand2_1
XFILLER_165_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19158_ _19158_/A _08947_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[28] sky130_fd_sc_hd__ebufn_8
XFILLER_34_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_1266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18109_ _18110_/CLK _18109_/D vssd1 vssd1 vccd1 vccd1 _18109_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_106_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_219_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_195_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_219_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_172_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09813_ _09813_/A _09813_/B vssd1 vssd1 vccd1 vccd1 _10366_/B sky130_fd_sc_hd__xnor2_2
XFILLER_143_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_228_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09744_ _09742_/A _09732_/B _09743_/X vssd1 vssd1 vccd1 vccd1 _09800_/B sky130_fd_sc_hd__a21o_1
XFILLER_132_1351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_228_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_215_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09675_ _18233_/Q _18232_/Q _18231_/Q vssd1 vssd1 vccd1 vccd1 _10600_/B sky130_fd_sc_hd__or3_4
XFILLER_55_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_227_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_230_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10450_ _09277_/A _09277_/B _10450_/S vssd1 vssd1 vccd1 vccd1 _10450_/X sky130_fd_sc_hd__mux2_1
XFILLER_202_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09109_ _09109_/A _09109_/B _09109_/C _09109_/D vssd1 vssd1 vccd1 vccd1 _09120_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_13_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10381_ _09309_/A _09319_/D _12124_/A vssd1 vssd1 vccd1 vccd1 _10381_/X sky130_fd_sc_hd__mux2_1
XFILLER_11_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12120_ _12120_/A _14267_/B vssd1 vssd1 vccd1 vccd1 _12120_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_163_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_190_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12051_ _12051_/A vssd1 vssd1 vccd1 vccd1 _13710_/A sky130_fd_sc_hd__buf_4
XFILLER_85_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11002_ _17822_/Q vssd1 vssd1 vccd1 vccd1 _11892_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_77_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19045__16 vssd1 vssd1 vccd1 vccd1 _19045__16/HI _19139_/A sky130_fd_sc_hd__conb_1
X_15810_ _15869_/A vssd1 vssd1 vccd1 vccd1 _15857_/A sky130_fd_sc_hd__clkbuf_2
X_16790_ _16792_/B _16788_/X _16789_/Y _16781_/X vssd1 vssd1 vccd1 vccd1 _18766_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_218_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15741_ _15743_/B _15737_/X _15738_/Y _15740_/X vssd1 vssd1 vccd1 vccd1 _18514_/D
+ sky130_fd_sc_hd__o211a_1
X_12953_ _12950_/Y _12935_/X _12951_/Y _17983_/Q _12952_/X vssd1 vssd1 vccd1 vccd1
+ _12953_/X sky130_fd_sc_hd__o221a_1
XTAP_3220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_219_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11904_ _11281_/B _11947_/B _12041_/B vssd1 vssd1 vccd1 vccd1 _11973_/A sky130_fd_sc_hd__o21ai_4
X_15672_ _18533_/Q _18497_/Q _15693_/S vssd1 vssd1 vccd1 vccd1 _15672_/X sky130_fd_sc_hd__mux2_1
X_18460_ _18467_/CLK _18460_/D vssd1 vssd1 vccd1 vccd1 _18460_/Q sky130_fd_sc_hd__dfxtp_2
Xclkbuf_leaf_42_wb_clk_i clkbuf_5_18_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18799_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_3264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12884_ _17958_/Q _12886_/C _12874_/X vssd1 vssd1 vccd1 vccd1 _12884_/Y sky130_fd_sc_hd__o21ai_1
XTAP_2530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14623_ _17687_/A _17663_/B vssd1 vssd1 vccd1 vccd1 _16886_/A sky130_fd_sc_hd__or2_4
XTAP_2563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17411_ _17472_/A vssd1 vssd1 vccd1 vccd1 _17538_/C sky130_fd_sc_hd__clkbuf_2
X_18391_ _18392_/CLK _18391_/D vssd1 vssd1 vccd1 vccd1 _18391_/Q sky130_fd_sc_hd__dfxtp_2
X_11835_ _11508_/C _11730_/B _11413_/Y _11834_/X _11828_/Y vssd1 vssd1 vccd1 vccd1
+ _11835_/X sky130_fd_sc_hd__a32o_1
XFILLER_2_1294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17342_ _17349_/B _17339_/X _17340_/X _17341_/X vssd1 vssd1 vccd1 vccd1 _18897_/D
+ sky130_fd_sc_hd__o211a_1
X_14554_ _16823_/A vssd1 vssd1 vccd1 vccd1 _15162_/B sky130_fd_sc_hd__buf_6
XFILLER_18_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11766_ _11757_/A _11797_/A _11763_/X _11765_/X vssd1 vssd1 vccd1 vccd1 _11766_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_53_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13505_ _13505_/A vssd1 vssd1 vccd1 vccd1 _13869_/A sky130_fd_sc_hd__buf_6
XFILLER_41_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10717_ _10781_/S vssd1 vssd1 vccd1 vccd1 _10883_/B sky130_fd_sc_hd__buf_4
X_17273_ _17273_/A _17275_/B vssd1 vssd1 vccd1 vccd1 _17273_/Y sky130_fd_sc_hd__nand2_1
XFILLER_202_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14485_ _18217_/Q _14491_/B vssd1 vssd1 vccd1 vccd1 _14486_/A sky130_fd_sc_hd__and2_1
X_11697_ _11696_/C _11685_/X _11687_/Y _11696_/X vssd1 vssd1 vccd1 vccd1 _11697_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_105_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16224_ _16356_/B vssd1 vssd1 vccd1 vccd1 _16272_/C sky130_fd_sc_hd__clkbuf_2
X_19012_ _19029_/CLK _19012_/D vssd1 vssd1 vccd1 vccd1 _19012_/Q sky130_fd_sc_hd__dfxtp_1
X_13436_ _13436_/A _13436_/B _13436_/C vssd1 vssd1 vccd1 vccd1 _13438_/C sky130_fd_sc_hd__or3_1
X_10648_ _10764_/A vssd1 vssd1 vccd1 vccd1 _10648_/X sky130_fd_sc_hd__buf_4
XFILLER_173_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16155_ _16160_/B _16152_/X _16154_/X _16139_/X vssd1 vssd1 vccd1 vccd1 _18612_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_173_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13367_ _13367_/A vssd1 vssd1 vccd1 vccd1 _17768_/A sky130_fd_sc_hd__clkbuf_2
X_10579_ _10572_/X _10578_/X _12061_/A vssd1 vssd1 vccd1 vccd1 _10579_/X sky130_fd_sc_hd__o21a_1
XFILLER_155_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15106_ _18401_/Q _18365_/Q _15121_/S vssd1 vssd1 vccd1 vccd1 _15106_/X sky130_fd_sc_hd__mux2_1
XFILLER_127_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12318_ _13037_/A vssd1 vssd1 vccd1 vccd1 _12318_/X sky130_fd_sc_hd__buf_6
X_16086_ _16689_/A _16150_/B vssd1 vssd1 vccd1 vccd1 _16096_/B sky130_fd_sc_hd__nor2_2
XFILLER_5_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13298_ _13298_/A _13298_/B vssd1 vssd1 vccd1 vccd1 _13311_/B sky130_fd_sc_hd__or2_1
XFILLER_114_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15037_ _18383_/Q _18347_/Q _15052_/S vssd1 vssd1 vccd1 vccd1 _15037_/X sky130_fd_sc_hd__mux2_1
X_12249_ _12249_/A vssd1 vssd1 vccd1 vccd1 _17861_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_29_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_229_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_231_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16988_ _18135_/Q _17278_/B vssd1 vssd1 vccd1 vccd1 _17098_/A sky130_fd_sc_hd__nand2_1
XFILLER_7_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18727_ _18738_/CLK _18727_/D vssd1 vssd1 vccd1 vccd1 _18727_/Q sky130_fd_sc_hd__dfxtp_1
X_15939_ _15942_/B _15937_/X _15938_/Y _15925_/X vssd1 vssd1 vccd1 vccd1 _18562_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_83_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_225_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09460_ _09475_/B vssd1 vssd1 vccd1 vccd1 _09461_/A sky130_fd_sc_hd__buf_2
XFILLER_224_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18658_ _18658_/CLK _18658_/D vssd1 vssd1 vccd1 vccd1 _18658_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_149_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_212_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17609_ _17567_/X _17602_/Y _17603_/X _17605_/Y _18964_/Q vssd1 vssd1 vccd1 vccd1
+ _17610_/B sky130_fd_sc_hd__a32o_1
XFILLER_224_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09391_ _18350_/Q _18349_/Q _18348_/Q vssd1 vssd1 vccd1 vccd1 _09392_/D sky130_fd_sc_hd__or3_4
XFILLER_149_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18589_ _18590_/CLK _18589_/D vssd1 vssd1 vccd1 vccd1 _18589_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_52_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_225_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_225_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_178_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_192_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_160_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_218_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_219_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_219_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_216_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09727_ _12063_/A _10033_/A vssd1 vssd1 vccd1 vccd1 _09728_/D sky130_fd_sc_hd__nor2_4
XFILLER_28_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09658_ _18109_/Q _17976_/Q vssd1 vssd1 vccd1 vccd1 _09659_/B sky130_fd_sc_hd__xnor2_1
XFILLER_227_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_216_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_215_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_231_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09589_ _10038_/B _09589_/B vssd1 vssd1 vccd1 vccd1 _09723_/A sky130_fd_sc_hd__and2b_4
XFILLER_163_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11620_ _11610_/Y _11618_/Y _11619_/X vssd1 vssd1 vccd1 vccd1 _11620_/Y sky130_fd_sc_hd__o21bai_1
XFILLER_179_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_211_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_196_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11551_ _17866_/Q vssd1 vssd1 vccd1 vccd1 _12267_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_204_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10502_ _10443_/X _10487_/X _10493_/X _10501_/X vssd1 vssd1 vccd1 vccd1 _10502_/X
+ sky130_fd_sc_hd__a211o_1
X_14270_ _14533_/A vssd1 vssd1 vccd1 vccd1 _14270_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_11482_ _11482_/A _11482_/B vssd1 vssd1 vccd1 vccd1 _11483_/C sky130_fd_sc_hd__nand2_1
XFILLER_10_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_160_wb_clk_i _18114_/CLK vssd1 vssd1 vccd1 vccd1 _17987_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_137_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13221_ _13221_/A vssd1 vssd1 vccd1 vccd1 _18065_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_136_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10433_ _10475_/A vssd1 vssd1 vccd1 vccd1 _10926_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_13_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13152_ _13152_/A vssd1 vssd1 vccd1 vccd1 _18034_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_109_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10364_ _10362_/X _10363_/X _10370_/S vssd1 vssd1 vccd1 vccd1 _10364_/X sky130_fd_sc_hd__mux2_1
XFILLER_174_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12103_ _12103_/A _12103_/B _12103_/C _12103_/D vssd1 vssd1 vccd1 vccd1 _12104_/D
+ sky130_fd_sc_hd__or4_1
XFILLER_174_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13083_ _13083_/A vssd1 vssd1 vccd1 vccd1 _18004_/D sky130_fd_sc_hd__clkbuf_1
X_17960_ _17965_/CLK _17960_/D vssd1 vssd1 vccd1 vccd1 _17960_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_88_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_215_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10295_ _09193_/A _09958_/A _10293_/X _10294_/X vssd1 vssd1 vccd1 vccd1 _10295_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_3_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16911_ _16916_/B _16908_/X _16910_/X _16893_/X vssd1 vssd1 vccd1 vccd1 _18792_/D
+ sky130_fd_sc_hd__o211a_1
X_12034_ _10236_/X _12092_/B _12012_/Y _12031_/Y _12033_/Y vssd1 vssd1 vccd1 vccd1
+ _12034_/X sky130_fd_sc_hd__a2111o_1
XFILLER_215_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17891_ _17891_/CLK _17891_/D vssd1 vssd1 vccd1 vccd1 _17891_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_2_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_211_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_215_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16842_ _18814_/Q _18778_/Q _16842_/S vssd1 vssd1 vccd1 vccd1 _16842_/X sky130_fd_sc_hd__mux2_1
XFILLER_78_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13985_ _18394_/Q _13522_/A _13630_/A _18376_/Q vssd1 vssd1 vccd1 vccd1 _13985_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_168_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16773_ _16796_/A _16773_/B _16773_/C vssd1 vssd1 vccd1 vccd1 _16773_/X sky130_fd_sc_hd__or3_1
X_18512_ _18548_/CLK _18512_/D vssd1 vssd1 vccd1 vccd1 _18512_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_111_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15724_ _15734_/A _16021_/B _15724_/C vssd1 vssd1 vccd1 vccd1 _15724_/X sky130_fd_sc_hd__or3_1
X_12936_ _17994_/Q _12955_/A vssd1 vssd1 vccd1 vccd1 _12936_/Y sky130_fd_sc_hd__nand2_1
XFILLER_59_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18443_ _18443_/CLK _18443_/D vssd1 vssd1 vccd1 vccd1 _18443_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_185_1366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15655_ _15678_/A _15946_/B _15666_/C vssd1 vssd1 vccd1 vccd1 _15655_/X sky130_fd_sc_hd__or3_1
XFILLER_209_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12867_ _12868_/B _12867_/B vssd1 vssd1 vccd1 vccd1 _17952_/D sky130_fd_sc_hd__nor2_1
XFILLER_61_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_222_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14606_ _14606_/A _14606_/B vssd1 vssd1 vccd1 vccd1 _14606_/Y sky130_fd_sc_hd__nand2_1
XFILLER_15_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11818_ _11742_/A _11742_/B _11742_/C vssd1 vssd1 vccd1 vccd1 _11818_/Y sky130_fd_sc_hd__o21ai_1
X_15586_ _18513_/Q _18477_/Q _15586_/S vssd1 vssd1 vccd1 vccd1 _15586_/X sky130_fd_sc_hd__mux2_1
X_18374_ _18374_/CLK _18374_/D vssd1 vssd1 vccd1 vccd1 _18374_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_1670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12798_ _17966_/Q vssd1 vssd1 vccd1 vccd1 _12798_/Y sky130_fd_sc_hd__inv_2
XFILLER_222_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14537_ _15643_/A vssd1 vssd1 vccd1 vccd1 _17541_/A sky130_fd_sc_hd__buf_2
XFILLER_18_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17325_ _17327_/B _17321_/X _17322_/Y _17324_/X vssd1 vssd1 vccd1 vccd1 _18892_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_230_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11749_ _11749_/A _11749_/B _11749_/C vssd1 vssd1 vccd1 vccd1 _11856_/B sky130_fd_sc_hd__nor3_1
XFILLER_187_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14468_ _14470_/B _14470_/C _14467_/Y vssd1 vssd1 vccd1 vccd1 _18209_/D sky130_fd_sc_hd__a21oi_1
X_17256_ _17256_/A _17538_/B _17256_/C vssd1 vssd1 vccd1 vccd1 _17256_/X sky130_fd_sc_hd__or3_1
XFILLER_146_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16207_ _16962_/A vssd1 vssd1 vccd1 vccd1 _16796_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_128_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13419_ _13415_/Y _13418_/X _18153_/Q _10990_/X vssd1 vssd1 vccd1 vccd1 _18153_/D
+ sky130_fd_sc_hd__a2bb2o_1
X_17187_ _17210_/A _17189_/B vssd1 vssd1 vccd1 vccd1 _17187_/Y sky130_fd_sc_hd__nand2_1
X_14399_ _14399_/A vssd1 vssd1 vccd1 vccd1 _14423_/A sky130_fd_sc_hd__clkbuf_2
X_16138_ _16181_/A _16736_/B _16181_/C vssd1 vssd1 vccd1 vccd1 _16138_/X sky130_fd_sc_hd__or3_1
XFILLER_142_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16069_ _16197_/A vssd1 vssd1 vccd1 vccd1 _16173_/A sky130_fd_sc_hd__clkbuf_2
X_08960_ _08960_/A vssd1 vssd1 vccd1 vccd1 _08960_/Y sky130_fd_sc_hd__inv_2
XFILLER_170_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09512_ _17591_/A vssd1 vssd1 vccd1 vccd1 _14386_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_225_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_224_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09443_ _09443_/A vssd1 vssd1 vccd1 vccd1 _09443_/Y sky130_fd_sc_hd__inv_2
XFILLER_64_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_213_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_212_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_225_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09374_ _18398_/Q _18397_/Q _18396_/Q vssd1 vssd1 vccd1 vccd1 _09376_/C sky130_fd_sc_hd__or3_4
XFILLER_75_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_203_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10080_ _09728_/D _10078_/X _10079_/X _10966_/B vssd1 vssd1 vccd1 vccd1 _10080_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_5914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_0 wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_5925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_181_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_1306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13770_ _18516_/Q _13759_/X _13732_/X _18507_/Q _13769_/X vssd1 vssd1 vccd1 vccd1
+ _13770_/X sky130_fd_sc_hd__a221o_2
X_10982_ _10982_/A vssd1 vssd1 vccd1 vccd1 _10982_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_90_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_231_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12721_ _12775_/A vssd1 vssd1 vccd1 vccd1 _12721_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_55_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_231_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15440_ _15440_/A vssd1 vssd1 vccd1 vccd1 _15458_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_203_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12652_ _17933_/Q _12653_/B vssd1 vssd1 vccd1 vccd1 _12654_/A sky130_fd_sc_hd__nor2_1
XFILLER_128_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11603_ _11603_/A _11603_/B vssd1 vssd1 vccd1 vccd1 _11603_/Y sky130_fd_sc_hd__nand2_1
X_15371_ _15423_/A _15371_/B _15423_/C vssd1 vssd1 vccd1 vccd1 _15371_/X sky130_fd_sc_hd__or3_1
XFILLER_212_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_208_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12583_ _12635_/A vssd1 vssd1 vccd1 vccd1 _12613_/A sky130_fd_sc_hd__buf_2
XFILLER_169_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_184_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17110_ _17115_/B _17108_/X _17109_/X _17096_/X vssd1 vssd1 vccd1 vccd1 _18840_/D
+ sky130_fd_sc_hd__o211a_1
X_14322_ _14334_/A _14322_/B vssd1 vssd1 vccd1 vccd1 _14322_/Y sky130_fd_sc_hd__nand2_1
XFILLER_211_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11534_ _11534_/A _11534_/B vssd1 vssd1 vccd1 vccd1 _11534_/Y sky130_fd_sc_hd__nor2_1
X_18090_ _18224_/CLK _18090_/D vssd1 vssd1 vccd1 vccd1 _18090_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_89_1307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17041_ _18822_/Q _17046_/B _17039_/X _17040_/X vssd1 vssd1 vccd1 vccd1 _18822_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_183_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14253_ _14203_/X _14249_/X _14305_/B _14219_/X vssd1 vssd1 vccd1 vccd1 _14253_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_125_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11465_ _11828_/A _11459_/X _11464_/X vssd1 vssd1 vccd1 vccd1 _11465_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_171_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13204_ _13208_/A _18059_/Q vssd1 vssd1 vccd1 vccd1 _13205_/A sky130_fd_sc_hd__and2_1
XFILLER_109_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10416_ _10555_/A vssd1 vssd1 vccd1 vccd1 _10932_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_171_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14184_ _18168_/Q _13409_/X _14113_/X _14183_/X vssd1 vssd1 vccd1 vccd1 _14185_/B
+ sky130_fd_sc_hd__o22ai_1
XFILLER_152_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11396_ _11595_/A _11396_/B vssd1 vssd1 vccd1 vccd1 _11730_/B sky130_fd_sc_hd__or2_4
XFILLER_180_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13135_ _13135_/A vssd1 vssd1 vccd1 vccd1 _18026_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_48_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10347_ _09114_/A _09109_/A _09119_/B _10728_/A _09923_/X _09935_/X vssd1 vssd1 vccd1
+ vccd1 _10347_/X sky130_fd_sc_hd__mux4_1
XTAP_706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18992_ _18992_/CLK _18992_/D vssd1 vssd1 vccd1 vccd1 _18992_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_79_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17943_ _18213_/CLK _17943_/D vssd1 vssd1 vccd1 vccd1 _17943_/Q sky130_fd_sc_hd__dfxtp_1
X_13066_ _13375_/A _13066_/B _13066_/C vssd1 vssd1 vccd1 vccd1 _13067_/A sky130_fd_sc_hd__and3_1
XFILLER_140_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10278_ _10278_/A vssd1 vssd1 vccd1 vccd1 _10278_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_97_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_1215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12017_ _12049_/A _12015_/Y _11999_/C _12016_/Y vssd1 vssd1 vccd1 vccd1 _12049_/B
+ sky130_fd_sc_hd__o2bb2a_2
XFILLER_152_1354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17874_ _19031_/CLK _17874_/D vssd1 vssd1 vccd1 vccd1 _17874_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_94_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_1338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16825_ _16871_/A vssd1 vssd1 vccd1 vccd1 _16825_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_120_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16756_ _16755_/B _16754_/X _16755_/Y _16740_/X vssd1 vssd1 vccd1 vccd1 _18758_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_59_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13968_ _18418_/Q _13651_/X _13964_/X _13967_/X vssd1 vssd1 vccd1 vccd1 _13968_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_222_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15707_ _15889_/A vssd1 vssd1 vccd1 vccd1 _15754_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_34_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12919_ _12987_/A _12919_/B vssd1 vssd1 vccd1 vccd1 _12919_/X sky130_fd_sc_hd__and2b_1
XFILLER_34_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13899_ _18541_/Q _13848_/A _13580_/A _18535_/Q _13898_/X vssd1 vssd1 vccd1 vccd1
+ _13899_/X sky130_fd_sc_hd__a221o_1
X_16687_ _16686_/B _16685_/X _16686_/Y _16683_/X vssd1 vssd1 vccd1 vccd1 _18740_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_146_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_222_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18426_ _18434_/CLK _18426_/D vssd1 vssd1 vccd1 vccd1 _18426_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_185_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15638_ _15678_/A _15935_/B _15666_/C vssd1 vssd1 vccd1 vccd1 _15638_/X sky130_fd_sc_hd__or3_1
XFILLER_21_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18357_ _18387_/CLK _18357_/D vssd1 vssd1 vccd1 vccd1 _18357_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_21_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15569_ _18509_/Q _18473_/Q _15586_/S vssd1 vssd1 vccd1 vccd1 _15569_/X sky130_fd_sc_hd__mux2_1
XFILLER_148_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17308_ _17318_/A _17449_/B _17318_/C vssd1 vssd1 vccd1 vccd1 _17308_/X sky130_fd_sc_hd__or3_1
XFILLER_174_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09090_ _18791_/Q _18790_/Q _18789_/Q vssd1 vssd1 vccd1 vccd1 _09093_/B sky130_fd_sc_hd__or3_4
XFILLER_148_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18288_ _18296_/CLK _18288_/D vssd1 vssd1 vccd1 vccd1 _18288_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_147_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17239_ _18908_/Q _18872_/Q _17244_/S vssd1 vssd1 vccd1 vccd1 _17239_/X sky130_fd_sc_hd__mux2_1
XFILLER_163_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09992_ _10103_/B vssd1 vssd1 vccd1 vccd1 _10004_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_143_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_192_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08943_ _08967_/A vssd1 vssd1 vccd1 vccd1 _08948_/A sky130_fd_sc_hd__buf_12
XFILLER_130_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_215_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_225_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09426_ _09482_/A vssd1 vssd1 vccd1 vccd1 _18146_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_52_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_212_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_198_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_212_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09357_ _18299_/Q _18298_/Q _18297_/Q vssd1 vssd1 vccd1 vccd1 _09360_/B sky130_fd_sc_hd__or3_2
XFILLER_205_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09288_ _09288_/A _09288_/B _09288_/C vssd1 vssd1 vccd1 vccd1 _09432_/C sky130_fd_sc_hd__nand3_2
XFILLER_14_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11250_ _11359_/B _11404_/B vssd1 vssd1 vccd1 vccd1 _11405_/A sky130_fd_sc_hd__or2_1
XFILLER_88_1351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10201_ _10201_/A _10201_/B vssd1 vssd1 vccd1 vccd1 _10202_/B sky130_fd_sc_hd__and2_1
XFILLER_175_1354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11181_ _11181_/A _11184_/C vssd1 vssd1 vccd1 vccd1 _11182_/C sky130_fd_sc_hd__or2_1
XFILLER_49_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_1207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10132_ _10456_/A _10441_/A _10131_/Y vssd1 vssd1 vccd1 vccd1 _10175_/A sky130_fd_sc_hd__a21o_2
XTAP_5700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14940_ _14975_/A _15233_/B _14965_/C vssd1 vssd1 vccd1 vccd1 _14940_/X sky130_fd_sc_hd__or3_1
X_10063_ _09160_/A _10040_/A _09999_/A _09193_/B _09688_/A vssd1 vssd1 vccd1 vccd1
+ _10063_/X sky130_fd_sc_hd__a221o_1
XFILLER_88_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14871_ _18343_/Q _18307_/Q _14883_/S vssd1 vssd1 vccd1 vccd1 _14871_/X sky130_fd_sc_hd__mux2_1
XTAP_5799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16610_ _18758_/Q _18722_/Q _16617_/S vssd1 vssd1 vccd1 vccd1 _16610_/X sky130_fd_sc_hd__mux2_1
XFILLER_63_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13822_ _18558_/Q _13735_/A _13764_/A _18582_/Q vssd1 vssd1 vccd1 vccd1 _13822_/X
+ sky130_fd_sc_hd__a22o_1
X_17590_ _17635_/A _17687_/B vssd1 vssd1 vccd1 vccd1 _17590_/Y sky130_fd_sc_hd__nor2_2
XFILLER_217_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_1322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_216_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_107 _13940_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16541_ _16578_/A vssd1 vssd1 vccd1 vccd1 _16602_/B sky130_fd_sc_hd__clkbuf_2
X_13753_ _18774_/Q _13719_/X _13752_/X _18780_/Q vssd1 vssd1 vccd1 vccd1 _13753_/X
+ sky130_fd_sc_hd__a22o_1
XINSDIODE2_118 _17471_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_129 _16219_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10965_ _09720_/X _10945_/X _10949_/X _10964_/X vssd1 vssd1 vccd1 vccd1 _10965_/Y
+ sky130_fd_sc_hd__a31oi_4
XFILLER_188_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12704_ _12698_/Y _12702_/X _12707_/C vssd1 vssd1 vccd1 vccd1 _12704_/X sky130_fd_sc_hd__o21ba_1
X_16472_ _16475_/B _16470_/X _16471_/Y _16456_/X vssd1 vssd1 vccd1 vccd1 _18688_/D
+ sky130_fd_sc_hd__o211a_1
X_13684_ _13684_/A vssd1 vssd1 vccd1 vccd1 _13684_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_188_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10896_ _10850_/X _10889_/X _10895_/X _12056_/A vssd1 vssd1 vccd1 vccd1 _10896_/Y
+ sky130_fd_sc_hd__a22oi_1
XFILLER_182_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18211_ _18213_/CLK _18211_/D vssd1 vssd1 vccd1 vccd1 _18211_/Q sky130_fd_sc_hd__dfxtp_1
X_15423_ _15423_/A _16021_/B _15423_/C vssd1 vssd1 vccd1 vccd1 _15423_/X sky130_fd_sc_hd__or3_1
X_12635_ _12635_/A vssd1 vssd1 vccd1 vccd1 _12635_/X sky130_fd_sc_hd__clkbuf_2
X_19191_ _19191_/A _08991_/Y vssd1 vssd1 vccd1 vccd1 io_out[29] sky130_fd_sc_hd__ebufn_8
XFILLER_12_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15354_ _16865_/A vssd1 vssd1 vccd1 vccd1 _15962_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_169_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18142_ _18147_/CLK _18142_/D vssd1 vssd1 vccd1 vccd1 _18142_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_180_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12566_ _12561_/Y _12563_/Y _12565_/X vssd1 vssd1 vccd1 vccd1 _12566_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_54_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_180_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11517_ _17871_/Q _17870_/Q vssd1 vssd1 vccd1 vccd1 _12285_/B sky130_fd_sc_hd__or2_1
X_14305_ _14305_/A _14305_/B vssd1 vssd1 vccd1 vccd1 _14305_/Y sky130_fd_sc_hd__nor2_1
XFILLER_102_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15285_ _18446_/Q _18410_/Q _15285_/S vssd1 vssd1 vccd1 vccd1 _15285_/X sky130_fd_sc_hd__mux2_1
XFILLER_144_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18073_ _18085_/CLK _18073_/D vssd1 vssd1 vccd1 vccd1 _18073_/Q sky130_fd_sc_hd__dfxtp_1
X_12497_ _12497_/A vssd1 vssd1 vccd1 vccd1 _17910_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_184_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_172_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17024_ _17023_/B _17022_/X _17023_/Y _17020_/X vssd1 vssd1 vccd1 vccd1 _18818_/D
+ sky130_fd_sc_hd__o211a_1
X_14236_ _18996_/Q _18998_/Q vssd1 vssd1 vccd1 vccd1 _14237_/A sky130_fd_sc_hd__nor2_1
XFILLER_144_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11448_ _11467_/D vssd1 vssd1 vccd1 vccd1 _11654_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_125_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14167_ _13710_/Y _14159_/X _14166_/X _13649_/X vssd1 vssd1 vccd1 vccd1 _14167_/X
+ sky130_fd_sc_hd__a22o_1
X_11379_ _11345_/A _17875_/Q _11331_/X _11329_/Y _11346_/Y vssd1 vssd1 vccd1 vccd1
+ _11379_/X sky130_fd_sc_hd__o311a_1
XFILLER_125_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13118_ _13118_/A _18020_/Q vssd1 vssd1 vccd1 vccd1 _13119_/A sky130_fd_sc_hd__and2_1
XTAP_514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14098_ _18644_/Q _13834_/A _13515_/A _18638_/Q _14097_/X vssd1 vssd1 vccd1 vccd1
+ _14098_/X sky130_fd_sc_hd__a221o_1
XFILLER_124_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18975_ _18977_/CLK _18975_/D vssd1 vssd1 vccd1 vccd1 _18975_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13049_ _13049_/A _13049_/B vssd1 vssd1 vccd1 vccd1 _13050_/A sky130_fd_sc_hd__and2_1
X_17926_ _17926_/CLK _17926_/D vssd1 vssd1 vccd1 vccd1 _17926_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_26_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17857_ _19034_/CLK _17857_/D vssd1 vssd1 vccd1 vccd1 _17857_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_187_1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16808_ _16808_/A vssd1 vssd1 vccd1 vccd1 _16866_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_82_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17788_ _17793_/CLK _17788_/D vssd1 vssd1 vccd1 vccd1 _17788_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_81_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_228_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16739_ _16752_/A _16743_/B vssd1 vssd1 vccd1 vccd1 _16739_/Y sky130_fd_sc_hd__nand2_1
XFILLER_81_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_223_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09211_ _18683_/Q _18682_/Q _18681_/Q vssd1 vssd1 vccd1 vccd1 _09214_/B sky130_fd_sc_hd__or3_4
X_18409_ _18443_/CLK _18409_/D vssd1 vssd1 vccd1 vccd1 _18409_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_14_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_194_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_179_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_222_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_195_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09142_ _18710_/Q _18709_/Q _18708_/Q vssd1 vssd1 vccd1 vccd1 _09143_/D sky130_fd_sc_hd__or3_4
XFILLER_135_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09073_ _09073_/A vssd1 vssd1 vccd1 vccd1 _19183_/A sky130_fd_sc_hd__buf_4
XFILLER_198_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_194_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_135_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09975_ _09969_/X _09971_/X _09973_/X _10356_/A vssd1 vssd1 vccd1 vccd1 _09975_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_226_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_217_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_213_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10750_ _10739_/X _10749_/X _10757_/B vssd1 vssd1 vccd1 vccd1 _10750_/X sky130_fd_sc_hd__mux2_1
XFILLER_213_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_198_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09409_ _18317_/Q _18316_/Q _18315_/Q vssd1 vssd1 vccd1 vccd1 _09413_/A sky130_fd_sc_hd__or3_2
XFILLER_55_1350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_185_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10681_ _09287_/A _09287_/D _09282_/D _09282_/B _10648_/X _12089_/A vssd1 vssd1 vccd1
+ vccd1 _10681_/X sky130_fd_sc_hd__mux4_2
XFILLER_164_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_139_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_199_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12420_ _17899_/Q _12420_/B _12420_/C vssd1 vssd1 vccd1 vccd1 _12420_/X sky130_fd_sc_hd__or3_1
XFILLER_205_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_224_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_205_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12351_ _12352_/B _12200_/X _12350_/Y vssd1 vssd1 vccd1 vccd1 _17891_/D sky130_fd_sc_hd__o21a_1
Xclkbuf_leaf_67_wb_clk_i clkbuf_5_20_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18708_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_181_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11302_ _11584_/B _11501_/A _11501_/C vssd1 vssd1 vccd1 vccd1 _11635_/A sky130_fd_sc_hd__or3_4
XFILLER_193_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15070_ _18355_/Q _15072_/B _15069_/Y _15066_/X vssd1 vssd1 vccd1 vccd1 _18355_/D
+ sky130_fd_sc_hd__o211a_1
X_12282_ _12282_/A vssd1 vssd1 vccd1 vccd1 _17870_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_135_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14021_ _18848_/Q _14019_/X _13842_/X _18854_/Q _14020_/X vssd1 vssd1 vccd1 vccd1
+ _14021_/X sky130_fd_sc_hd__a221o_1
XFILLER_4_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11233_ _11232_/B _11231_/A _11221_/X vssd1 vssd1 vccd1 vccd1 _11234_/B sky130_fd_sc_hd__o21ai_1
XFILLER_88_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_136_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11164_ _17816_/Q _17815_/Q _11164_/C _11164_/D vssd1 vssd1 vccd1 vccd1 _11212_/B
+ sky130_fd_sc_hd__nor4_4
XFILLER_136_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10115_ _10122_/A _10122_/B vssd1 vssd1 vccd1 vccd1 _10120_/B sky130_fd_sc_hd__or2_1
X_18760_ _18778_/CLK _18760_/D vssd1 vssd1 vccd1 vccd1 _18760_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_96_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15972_ _16028_/A vssd1 vssd1 vccd1 vccd1 _15972_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_5530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11095_ _12041_/A _11892_/B _11113_/S vssd1 vssd1 vccd1 vccd1 _11096_/A sky130_fd_sc_hd__mux2_1
XTAP_5541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17711_ _12972_/X _12770_/Y _12862_/X vssd1 vssd1 vccd1 vccd1 _18993_/D sky130_fd_sc_hd__a21oi_1
XFILLER_49_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14923_ _18319_/Q _14924_/B _14921_/Y _14922_/X vssd1 vssd1 vccd1 vccd1 _18319_/D
+ sky130_fd_sc_hd__o211a_1
X_10046_ _10046_/A vssd1 vssd1 vccd1 vccd1 _10090_/S sky130_fd_sc_hd__buf_4
XFILLER_76_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18691_ _18693_/CLK _18691_/D vssd1 vssd1 vccd1 vccd1 _18691_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_48_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17642_ _17641_/X _17635_/Y _17631_/X _17636_/Y _18973_/Q vssd1 vssd1 vccd1 vccd1
+ _17643_/B sky130_fd_sc_hd__a32o_1
XTAP_4873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14854_ _14918_/A vssd1 vssd1 vccd1 vccd1 _14985_/B sky130_fd_sc_hd__buf_2
XTAP_4884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_223_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_205_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13805_ _18390_/Q _13715_/A _13752_/A _18384_/Q vssd1 vssd1 vccd1 vccd1 _13805_/X
+ sky130_fd_sc_hd__a22o_1
X_17573_ _17587_/A _17573_/B vssd1 vssd1 vccd1 vccd1 _17574_/A sky130_fd_sc_hd__and2_1
X_14785_ _14810_/A _14788_/B vssd1 vssd1 vccd1 vccd1 _14785_/Y sky130_fd_sc_hd__nand2_1
X_11997_ _11997_/A _11999_/B vssd1 vssd1 vccd1 vccd1 _11997_/Y sky130_fd_sc_hd__nor2_1
XFILLER_95_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16524_ _16524_/A vssd1 vssd1 vccd1 vccd1 _16575_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_189_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13736_ _18318_/Q _13579_/A _13735_/X _18306_/Q vssd1 vssd1 vccd1 vccd1 _13736_/X
+ sky130_fd_sc_hd__a22o_1
X_10948_ _09408_/A _09408_/B _10948_/S vssd1 vssd1 vccd1 vccd1 _10948_/X sky130_fd_sc_hd__mux2_1
XFILLER_17_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_220_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16455_ _16491_/A _16749_/B _16481_/C vssd1 vssd1 vccd1 vccd1 _16455_/X sky130_fd_sc_hd__or3_1
XFILLER_188_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_177_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10879_ _10859_/S _10876_/X _10878_/X _10700_/S vssd1 vssd1 vccd1 vccd1 _10879_/X
+ sky130_fd_sc_hd__a211o_1
X_13667_ _13667_/A vssd1 vssd1 vccd1 vccd1 _13752_/A sky130_fd_sc_hd__buf_6
XFILLER_108_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15406_ _16922_/A vssd1 vssd1 vccd1 vccd1 _16005_/A sky130_fd_sc_hd__clkbuf_4
XPHY_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19174_ _19174_/A _09022_/Y vssd1 vssd1 vccd1 vccd1 io_out[12] sky130_fd_sc_hd__ebufn_8
X_12618_ _12618_/A _12618_/B vssd1 vssd1 vccd1 vccd1 _12619_/B sky130_fd_sc_hd__or2_1
X_16386_ _16434_/A _16678_/B _16422_/C vssd1 vssd1 vccd1 vccd1 _16386_/X sky130_fd_sc_hd__or3_1
XPHY_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13598_ _13630_/A vssd1 vssd1 vccd1 vccd1 _13598_/X sky130_fd_sc_hd__buf_6
XFILLER_118_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18125_ _18125_/CLK _18125_/D vssd1 vssd1 vccd1 vccd1 _18125_/Q sky130_fd_sc_hd__dfxtp_2
X_15337_ _15415_/A vssd1 vssd1 vccd1 vccd1 _15356_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_200_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12549_ _12542_/B _12523_/X _12545_/X _12547_/Y _12548_/X vssd1 vssd1 vccd1 vccd1
+ _17918_/D sky130_fd_sc_hd__a221o_1
XFILLER_144_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18056_ _18068_/CLK _18056_/D vssd1 vssd1 vccd1 vccd1 _18056_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_6_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15268_ _15279_/A _15268_/B _15279_/C vssd1 vssd1 vccd1 vccd1 _15268_/X sky130_fd_sc_hd__or3_1
XFILLER_144_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17007_ _17010_/B _17005_/X _17006_/Y _16999_/X vssd1 vssd1 vccd1 vccd1 _18814_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_6_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14219_ _14297_/A _14335_/B vssd1 vssd1 vccd1 vccd1 _14219_/X sky130_fd_sc_hd__and2_1
X_15199_ _15220_/A _15199_/B _15199_/C vssd1 vssd1 vccd1 vccd1 _15199_/X sky130_fd_sc_hd__or3_1
XFILLER_28_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_113_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09760_ _09760_/A _09760_/B vssd1 vssd1 vccd1 vccd1 _09760_/X sky130_fd_sc_hd__or2_1
XFILLER_101_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18958_ _18960_/CLK _18958_/D vssd1 vssd1 vccd1 vccd1 _18958_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_39_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17909_ _19034_/CLK _17909_/D vssd1 vssd1 vccd1 vccd1 _17909_/Q sky130_fd_sc_hd__dfxtp_1
X_09691_ _12068_/A _09691_/B vssd1 vssd1 vccd1 vccd1 _09691_/X sky130_fd_sc_hd__or2_1
X_18889_ _18893_/CLK _18889_/D vssd1 vssd1 vccd1 vccd1 _18889_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_94_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_215_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_215_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_212_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_176_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_148_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09125_ _18818_/Q _18817_/Q _18816_/Q vssd1 vssd1 vccd1 vccd1 _09126_/D sky130_fd_sc_hd__or3_4
XFILLER_157_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_198_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_159_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09056_ _09058_/A vssd1 vssd1 vccd1 vccd1 _09056_/Y sky130_fd_sc_hd__inv_2
XFILLER_136_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09958_ _09958_/A vssd1 vssd1 vccd1 vccd1 _10285_/S sky130_fd_sc_hd__buf_4
Xclkbuf_leaf_185_wb_clk_i clkbuf_5_8_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _19029_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_4103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_213_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_218_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_114_wb_clk_i clkbuf_5_31_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18458_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_09889_ _09889_/A vssd1 vssd1 vccd1 vccd1 _09889_/X sky130_fd_sc_hd__buf_2
XTAP_3402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11920_ _12120_/A _11920_/B vssd1 vssd1 vccd1 vccd1 _11920_/Y sky130_fd_sc_hd__nor2_1
XTAP_3435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11851_ _11598_/B _11683_/X _11829_/X _11859_/A _11850_/X vssd1 vssd1 vccd1 vccd1
+ _11851_/X sky130_fd_sc_hd__o311a_2
XFILLER_17_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10802_ _10805_/B _10801_/X _10818_/B vssd1 vssd1 vccd1 vccd1 _10802_/X sky130_fd_sc_hd__a21o_1
X_14570_ _14584_/A _14584_/B _15175_/B vssd1 vssd1 vccd1 vccd1 _14570_/X sky130_fd_sc_hd__or3_1
XFILLER_54_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11782_ _11770_/A _11784_/B _11770_/B vssd1 vssd1 vccd1 vccd1 _11783_/B sky130_fd_sc_hd__a21oi_1
XFILLER_220_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_213_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_201_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13521_ _13594_/A vssd1 vssd1 vccd1 vccd1 _13522_/A sky130_fd_sc_hd__buf_6
X_10733_ _10733_/A vssd1 vssd1 vccd1 vccd1 _10733_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_41_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_185_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16240_ _16265_/A _16243_/B vssd1 vssd1 vccd1 vccd1 _16240_/Y sky130_fd_sc_hd__nand2_1
X_13452_ _13452_/A _13452_/B vssd1 vssd1 vccd1 vccd1 _13452_/Y sky130_fd_sc_hd__nand2_1
XFILLER_9_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10664_ _10664_/A vssd1 vssd1 vccd1 vccd1 _10859_/S sky130_fd_sc_hd__buf_2
XFILLER_139_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_186_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12403_ _17897_/Q _12409_/B _12403_/C vssd1 vssd1 vccd1 vccd1 _12404_/B sky130_fd_sc_hd__nor3_1
XFILLER_90_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16171_ _16199_/A _16175_/B vssd1 vssd1 vccd1 vccd1 _16171_/Y sky130_fd_sc_hd__nand2_1
XFILLER_154_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13383_ _13383_/A vssd1 vssd1 vccd1 vccd1 _13383_/X sky130_fd_sc_hd__buf_2
X_10595_ _12063_/A _14317_/B vssd1 vssd1 vccd1 vccd1 _10595_/X sky130_fd_sc_hd__and2b_1
XFILLER_103_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_220_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15122_ _15162_/A _15268_/B _15136_/C vssd1 vssd1 vccd1 vccd1 _15122_/X sky130_fd_sc_hd__or3_1
X_12334_ _12334_/A vssd1 vssd1 vccd1 vccd1 _17884_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_86_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15053_ _15232_/A vssd1 vssd1 vccd1 vccd1 _15098_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_114_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12265_ _11563_/B _12261_/A _12261_/B vssd1 vssd1 vccd1 vccd1 _12270_/B sky130_fd_sc_hd__a21oi_1
XFILLER_147_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14004_ _18934_/Q _13785_/X _14002_/X _14003_/X vssd1 vssd1 vccd1 vccd1 _14004_/X
+ sky130_fd_sc_hd__a211o_1
X_11216_ _12361_/A vssd1 vssd1 vccd1 vccd1 _16891_/A sky130_fd_sc_hd__buf_12
X_12196_ _17906_/Q _17905_/Q _17904_/Q _17903_/Q vssd1 vssd1 vccd1 vccd1 _12476_/B
+ sky130_fd_sc_hd__or4_1
XFILLER_122_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18812_ _18812_/CLK _18812_/D vssd1 vssd1 vccd1 vccd1 _18812_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_6050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11147_ _11784_/A vssd1 vssd1 vccd1 vccd1 _11770_/A sky130_fd_sc_hd__buf_2
XTAP_6061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_228_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_1260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_163_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18743_ _18743_/CLK _18743_/D vssd1 vssd1 vccd1 vccd1 _18743_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15955_ _15960_/B _15950_/X _15954_/Y _15948_/X vssd1 vssd1 vccd1 vccd1 _18565_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_5360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11078_ _11078_/A vssd1 vssd1 vccd1 vccd1 _17789_/D sky130_fd_sc_hd__clkbuf_1
XTAP_5371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14906_ _14919_/A _15199_/B _14906_/C vssd1 vssd1 vccd1 vccd1 _14906_/X sky130_fd_sc_hd__or3_1
X_10029_ _10026_/X _10027_/X _10029_/S vssd1 vssd1 vccd1 vccd1 _10029_/X sky130_fd_sc_hd__mux2_1
XFILLER_76_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18674_ _18677_/CLK _18674_/D vssd1 vssd1 vccd1 vccd1 _18674_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_97_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_188_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15886_ _15938_/A _15890_/B vssd1 vssd1 vccd1 vccd1 _15886_/Y sky130_fd_sc_hd__nand2_1
XTAP_4670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17625_ _17575_/X _17623_/Y _17603_/X _17624_/Y _18969_/Q vssd1 vssd1 vccd1 vccd1
+ _17626_/B sky130_fd_sc_hd__a32o_1
XFILLER_184_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14837_ _18335_/Q _18299_/Q _14848_/S vssd1 vssd1 vccd1 vccd1 _14837_/X sky130_fd_sc_hd__mux2_1
XFILLER_63_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_184_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17556_ _17556_/A vssd1 vssd1 vccd1 vccd1 _17556_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_91_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14768_ _14767_/B _14765_/X _14767_/Y _14758_/X vssd1 vssd1 vccd1 vccd1 _18281_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_51_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_225_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16507_ _16507_/A _16510_/B vssd1 vssd1 vccd1 vccd1 _16507_/Y sky130_fd_sc_hd__nand2_1
XFILLER_16_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13719_ _13719_/A vssd1 vssd1 vccd1 vccd1 _13719_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_32_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17487_ _17489_/B _17485_/X _17486_/Y _17478_/X vssd1 vssd1 vccd1 vccd1 _18934_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_204_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14699_ _14948_/A vssd1 vssd1 vccd1 vccd1 _14753_/A sky130_fd_sc_hd__buf_4
XFILLER_225_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19226_ _19226_/A _08935_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[26] sky130_fd_sc_hd__ebufn_8
XFILLER_20_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16438_ _18679_/Q _16439_/B _16436_/Y _16437_/X vssd1 vssd1 vccd1 vccd1 _18679_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_149_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_1280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_220_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19157_ _19157_/A _08952_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[27] sky130_fd_sc_hd__ebufn_8
XFILLER_191_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16369_ _16433_/A vssd1 vssd1 vccd1 vccd1 _16501_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_157_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18108_ _18108_/CLK _18108_/D vssd1 vssd1 vccd1 vccd1 _18108_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_191_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_1327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18039_ _18094_/CLK _18039_/D vssd1 vssd1 vccd1 vccd1 _18039_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_114_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09812_ _09812_/A _09812_/B vssd1 vssd1 vccd1 vccd1 _09813_/B sky130_fd_sc_hd__xnor2_1
XFILLER_87_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_140_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_228_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09743_ _09743_/A _10705_/A vssd1 vssd1 vccd1 vccd1 _09743_/X sky130_fd_sc_hd__and2_1
XFILLER_132_1363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09674_ _10962_/A vssd1 vssd1 vccd1 vccd1 _12068_/A sky130_fd_sc_hd__buf_4
XFILLER_223_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_199_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_230_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_196_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_204_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09108_ _18770_/Q _18769_/Q _18768_/Q vssd1 vssd1 vccd1 vccd1 _09109_/D sky130_fd_sc_hd__or3_4
XFILLER_136_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10380_ _12126_/A _10374_/X _10378_/X _09889_/A _10379_/X vssd1 vssd1 vccd1 vccd1
+ _10380_/X sky130_fd_sc_hd__a32o_1
XFILLER_202_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09039_ _09040_/A vssd1 vssd1 vccd1 vccd1 _09039_/Y sky130_fd_sc_hd__inv_2
XFILLER_164_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12050_ _12055_/A _12055_/B _12055_/C _12055_/D vssd1 vssd1 vccd1 vccd1 _12051_/A
+ sky130_fd_sc_hd__or4_1
XFILLER_137_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11001_ _17819_/Q _11232_/B _11001_/C vssd1 vssd1 vccd1 vccd1 _11237_/B sky130_fd_sc_hd__and3_1
XFILLER_133_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_218_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15740_ _15823_/A vssd1 vssd1 vccd1 vccd1 _15740_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_3210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12952_ _12760_/A _12947_/X _12948_/X _12928_/X vssd1 vssd1 vccd1 vccd1 _12952_/X
+ sky130_fd_sc_hd__o31a_2
XFILLER_92_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11903_ _11947_/A vssd1 vssd1 vccd1 vccd1 _12041_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_93_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15671_ _15673_/B _15669_/X _15670_/Y _15662_/X vssd1 vssd1 vccd1 vccd1 _18496_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_3265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12883_ _12886_/C _12883_/B vssd1 vssd1 vccd1 vccd1 _17957_/D sky130_fd_sc_hd__nor2_1
XFILLER_73_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17410_ _17410_/A _17549_/B vssd1 vssd1 vccd1 vccd1 _17472_/A sky130_fd_sc_hd__or2_1
XTAP_3298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14622_ _14660_/B vssd1 vssd1 vccd1 vccd1 _17663_/B sky130_fd_sc_hd__clkbuf_2
XTAP_2553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18390_ _18392_/CLK _18390_/D vssd1 vssd1 vccd1 vccd1 _18390_/Q sky130_fd_sc_hd__dfxtp_2
X_11834_ _11582_/A _11396_/B _11413_/Y _11443_/X vssd1 vssd1 vccd1 vccd1 _11834_/X
+ sky130_fd_sc_hd__a31o_1
XTAP_2564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17341_ _17400_/A vssd1 vssd1 vccd1 vccd1 _17341_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_92_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14553_ _16817_/A vssd1 vssd1 vccd1 vccd1 _16823_/A sky130_fd_sc_hd__buf_6
X_11765_ _11261_/X _11730_/B _11764_/Y vssd1 vssd1 vccd1 vccd1 _11765_/X sky130_fd_sc_hd__o21a_1
Xclkbuf_leaf_82_wb_clk_i clkbuf_5_23_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18577_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_187_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13504_ _13719_/A vssd1 vssd1 vccd1 vccd1 _13505_/A sky130_fd_sc_hd__clkbuf_4
X_10716_ _10716_/A vssd1 vssd1 vccd1 vccd1 _10781_/S sky130_fd_sc_hd__buf_2
X_17272_ _18879_/Q _17275_/B _17271_/X _17260_/X vssd1 vssd1 vccd1 vccd1 _18879_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_159_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11696_ _11685_/X _11696_/B _11696_/C vssd1 vssd1 vccd1 vccd1 _11696_/X sky130_fd_sc_hd__and3b_1
X_14484_ _14484_/A vssd1 vssd1 vccd1 vccd1 _18216_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_11_wb_clk_i _17929_/CLK vssd1 vssd1 vccd1 vccd1 _17959_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_158_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19011_ _19029_/CLK _19011_/D vssd1 vssd1 vccd1 vccd1 _19011_/Q sky130_fd_sc_hd__dfxtp_1
X_16223_ _16289_/A vssd1 vssd1 vccd1 vccd1 _16356_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_173_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10647_ _10668_/A vssd1 vssd1 vccd1 vccd1 _10764_/A sky130_fd_sc_hd__buf_4
XFILLER_9_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13435_ _13710_/B _13435_/B vssd1 vssd1 vccd1 vccd1 _13436_/C sky130_fd_sc_hd__nor2_1
XFILLER_139_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_228_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16154_ _16181_/A _16749_/B _16181_/C vssd1 vssd1 vccd1 vccd1 _16154_/X sky130_fd_sc_hd__or3_1
XFILLER_6_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13366_ _18107_/Q _13336_/X _13370_/B vssd1 vssd1 vccd1 vccd1 _18107_/D sky130_fd_sc_hd__o21a_1
XFILLER_177_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10578_ _10029_/S _10573_/X _10577_/X _10009_/A vssd1 vssd1 vccd1 vccd1 _10578_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_127_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_182_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15105_ _15105_/A vssd1 vssd1 vccd1 vccd1 _15121_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_154_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12317_ _17879_/Q _11346_/A _12301_/A _12316_/X vssd1 vssd1 vccd1 vccd1 _12317_/Y
+ sky130_fd_sc_hd__o211ai_1
X_16085_ _16127_/A vssd1 vssd1 vccd1 vccd1 _16150_/B sky130_fd_sc_hd__buf_2
XFILLER_177_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13297_ _13297_/A _13297_/B _13297_/C vssd1 vssd1 vccd1 vccd1 _13298_/B sky130_fd_sc_hd__or3_1
XFILLER_5_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15036_ _15105_/A vssd1 vssd1 vccd1 vccd1 _15052_/S sky130_fd_sc_hd__clkbuf_2
X_12248_ _12517_/A _12248_/B vssd1 vssd1 vccd1 vccd1 _12249_/A sky130_fd_sc_hd__and2_1
XFILLER_64_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12179_ _12165_/Y _12175_/Y _12177_/X _12178_/X vssd1 vssd1 vccd1 vccd1 _17847_/D
+ sky130_fd_sc_hd__o31a_1
XFILLER_95_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_228_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16987_ _17423_/A _17109_/C vssd1 vssd1 vccd1 vccd1 _16998_/B sky130_fd_sc_hd__nor2_2
XFILLER_7_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_231_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18726_ _18738_/CLK _18726_/D vssd1 vssd1 vccd1 vccd1 _18726_/Q sky130_fd_sc_hd__dfxtp_1
X_15938_ _15938_/A _15942_/B vssd1 vssd1 vccd1 vccd1 _15938_/Y sky130_fd_sc_hd__nand2_1
XTAP_5190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_224_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18657_ _18663_/CLK _18657_/D vssd1 vssd1 vccd1 vccd1 _18657_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_92_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_225_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15869_ _15869_/A vssd1 vssd1 vccd1 vccd1 _15921_/A sky130_fd_sc_hd__buf_2
XFILLER_24_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_224_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_225_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17608_ _17608_/A vssd1 vssd1 vccd1 vccd1 _18963_/D sky130_fd_sc_hd__clkbuf_1
X_09390_ _18362_/Q _18361_/Q _18360_/Q vssd1 vssd1 vccd1 vccd1 _09392_/C sky130_fd_sc_hd__or3_2
XFILLER_24_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_212_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18588_ _18590_/CLK _18588_/D vssd1 vssd1 vccd1 vccd1 _18588_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_145_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_224_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17539_ _17544_/B _17537_/X _17538_/X _11816_/X vssd1 vssd1 vccd1 vccd1 _18948_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_225_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_1323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_225_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_1367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_178_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_220_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19209_ _19209_/A _08978_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[9] sky130_fd_sc_hd__ebufn_8
XFILLER_193_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_191_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_228_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09726_ _09726_/A _09726_/B vssd1 vssd1 vccd1 vccd1 _10033_/A sky130_fd_sc_hd__xnor2_4
XFILLER_216_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_227_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09657_ _09657_/A vssd1 vssd1 vccd1 vccd1 _09657_/X sky130_fd_sc_hd__buf_4
XFILLER_82_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09588_ _09725_/A _09725_/B vssd1 vssd1 vccd1 vccd1 _09588_/X sky130_fd_sc_hd__or2b_1
XTAP_1137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_169_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_208_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_179_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_168_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_196_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11550_ _17868_/Q vssd1 vssd1 vccd1 vccd1 _11565_/B sky130_fd_sc_hd__inv_2
XFILLER_184_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10501_ _10918_/S _10499_/X _10500_/X _10419_/A vssd1 vssd1 vccd1 vccd1 _10501_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_211_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_168_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11481_ _11318_/A _11477_/X _11480_/X _17888_/Q vssd1 vssd1 vccd1 vccd1 _11484_/A
+ sky130_fd_sc_hd__a211o_1
XFILLER_17_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_1240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13220_ _13222_/A _18066_/Q vssd1 vssd1 vccd1 vccd1 _13221_/A sky130_fd_sc_hd__and2_1
XFILLER_10_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10432_ _09136_/A _09126_/B _09131_/C _09136_/C _10429_/X _10430_/X vssd1 vssd1 vccd1
+ vccd1 _10432_/X sky130_fd_sc_hd__mux4_1
XFILLER_13_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13151_ _13151_/A _18035_/Q vssd1 vssd1 vccd1 vccd1 _13152_/A sky130_fd_sc_hd__and2_1
XFILLER_174_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10363_ _09103_/A _09098_/D _09093_/D _09103_/C _09953_/A _10375_/S vssd1 vssd1 vccd1
+ vccd1 _10363_/X sky130_fd_sc_hd__mux4_1
XFILLER_151_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19105__76 vssd1 vssd1 vccd1 vccd1 _19105__76/HI _19213_/A sky130_fd_sc_hd__conb_1
X_12102_ _12102_/A _12102_/B vssd1 vssd1 vccd1 vccd1 _12103_/D sky130_fd_sc_hd__xnor2_1
XFILLER_151_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_139_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13082_ _13082_/A _17517_/A vssd1 vssd1 vccd1 vccd1 _13083_/A sky130_fd_sc_hd__and2_1
XFILLER_151_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10294_ _10294_/A vssd1 vssd1 vccd1 vccd1 _10294_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_215_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16910_ _16936_/A _17493_/B _16936_/C vssd1 vssd1 vccd1 vccd1 _16910_/X sky130_fd_sc_hd__or3_1
XFILLER_2_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12033_ _10236_/X _12092_/B _12032_/X vssd1 vssd1 vccd1 vccd1 _12033_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_105_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17890_ _17890_/CLK _17890_/D vssd1 vssd1 vccd1 vccd1 _17890_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_78_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_215_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16841_ _16847_/B _16838_/X _16840_/X _16825_/X vssd1 vssd1 vccd1 vccd1 _18777_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_144_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16772_ _18798_/Q _18762_/Q _16784_/S vssd1 vssd1 vccd1 vccd1 _16772_/X sky130_fd_sc_hd__mux2_1
XFILLER_225_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13984_ _18370_/Q _13940_/A _13730_/A _18373_/Q _13983_/X vssd1 vssd1 vccd1 vccd1
+ _13984_/X sky130_fd_sc_hd__a221o_1
XFILLER_4_1346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18511_ _18511_/CLK _18511_/D vssd1 vssd1 vccd1 vccd1 _18511_/Q sky130_fd_sc_hd__dfxtp_2
X_15723_ _18546_/Q _18510_/Q _15733_/S vssd1 vssd1 vccd1 vccd1 _15723_/X sky130_fd_sc_hd__mux2_1
XFILLER_185_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12935_ _12951_/A vssd1 vssd1 vccd1 vccd1 _12935_/X sky130_fd_sc_hd__buf_2
XFILLER_80_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_1266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18442_ _18448_/CLK _18442_/D vssd1 vssd1 vccd1 vccd1 _18442_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_46_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15654_ _18528_/Q _18492_/Q _15665_/S vssd1 vssd1 vccd1 vccd1 _15654_/X sky130_fd_sc_hd__mux2_1
XFILLER_179_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12866_ _17952_/Q _12864_/A _12862_/X vssd1 vssd1 vccd1 vccd1 _12867_/B sky130_fd_sc_hd__o21ai_1
XTAP_2361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14605_ _18244_/Q _14606_/B _14604_/Y _14587_/X vssd1 vssd1 vccd1 vccd1 _18244_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_18_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18373_ _18373_/CLK _18373_/D vssd1 vssd1 vccd1 vccd1 _18373_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_21_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11817_ _11717_/Y _11810_/X _11813_/Y _18154_/Q _11816_/X vssd1 vssd1 vccd1 vccd1
+ _17825_/D sky130_fd_sc_hd__o221a_1
XTAP_2394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15585_ _16030_/A _15597_/B vssd1 vssd1 vccd1 vccd1 _15594_/B sky130_fd_sc_hd__nor2_2
XTAP_1660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12797_ _12676_/B _12795_/Y _12796_/Y _17935_/Q _17969_/Q vssd1 vssd1 vccd1 vccd1
+ _12797_/X sky130_fd_sc_hd__a221o_1
XTAP_1682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17324_ _17400_/A vssd1 vssd1 vccd1 vccd1 _17324_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_222_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14536_ _15951_/A vssd1 vssd1 vccd1 vccd1 _15643_/A sky130_fd_sc_hd__buf_12
XTAP_1693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11748_ _13446_/A _11748_/B _11748_/C vssd1 vssd1 vccd1 vccd1 _11749_/C sky130_fd_sc_hd__and3_1
XFILLER_230_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17255_ _18912_/Q _18876_/Q _17262_/S vssd1 vssd1 vccd1 vccd1 _17255_/X sky130_fd_sc_hd__mux2_1
XFILLER_179_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14467_ _14470_/B _14470_/C _14436_/A vssd1 vssd1 vccd1 vccd1 _14467_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_70_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11679_ _11664_/X _11677_/X _11845_/A vssd1 vssd1 vccd1 vccd1 _11680_/D sky130_fd_sc_hd__a21oi_1
X_16206_ _18660_/Q _18624_/Q _16215_/S vssd1 vssd1 vccd1 vccd1 _16206_/X sky130_fd_sc_hd__mux2_1
XFILLER_31_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13418_ _14355_/B _13418_/B _13418_/C _13418_/D vssd1 vssd1 vccd1 vccd1 _13418_/X
+ sky130_fd_sc_hd__or4_1
XFILLER_190_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17186_ _18858_/Q _17189_/B _17185_/X _17181_/X vssd1 vssd1 vccd1 vccd1 _18858_/D
+ sky130_fd_sc_hd__o211a_1
X_14398_ _14414_/A _14391_/Y _14386_/B vssd1 vssd1 vccd1 vccd1 _14398_/Y sky130_fd_sc_hd__o21bai_1
Xclkbuf_leaf_217_wb_clk_i clkbuf_5_8_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _19030_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_16137_ _16889_/A vssd1 vssd1 vccd1 vccd1 _16736_/B sky130_fd_sc_hd__buf_4
XFILLER_31_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13349_ _13346_/X _13348_/Y _17768_/B vssd1 vssd1 vccd1 vccd1 _18100_/D sky130_fd_sc_hd__a21boi_1
XFILLER_115_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16068_ _18141_/Q _16528_/B vssd1 vssd1 vccd1 vccd1 _16197_/A sky130_fd_sc_hd__nand2_1
XFILLER_103_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15019_ _15042_/A _15162_/B _15054_/C vssd1 vssd1 vccd1 vccd1 _15019_/X sky130_fd_sc_hd__or3_1
XFILLER_25_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_229_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_216_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09511_ _12217_/A vssd1 vssd1 vccd1 vccd1 _12257_/A sky130_fd_sc_hd__buf_2
X_18709_ _18710_/CLK _18709_/D vssd1 vssd1 vccd1 vccd1 _18709_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_204_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_225_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09442_ _09294_/X _09299_/X _09304_/X _09321_/A vssd1 vssd1 vccd1 vccd1 _09442_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_52_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_224_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_220_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09373_ _18383_/Q _18382_/Q _18381_/Q vssd1 vssd1 vccd1 vccd1 _09376_/B sky130_fd_sc_hd__or3_4
XFILLER_224_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_220_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_149_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_181_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_1 _16880_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_114_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_1318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_216_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09709_ _09709_/A vssd1 vssd1 vccd1 vccd1 _09709_/X sky130_fd_sc_hd__buf_4
XFILLER_62_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10981_ _14272_/A _15840_/A _14272_/B vssd1 vssd1 vccd1 vccd1 _10982_/A sky130_fd_sc_hd__and3_1
XFILLER_114_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12720_ _12926_/A vssd1 vssd1 vccd1 vccd1 _12775_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_71_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_231_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_204_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_216_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12651_ _12646_/B _12635_/X _12649_/Y _12650_/X _12621_/X vssd1 vssd1 vccd1 vccd1
+ _17929_/D sky130_fd_sc_hd__a221o_1
XFILLER_231_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_1340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11602_ _11615_/A _11602_/B vssd1 vssd1 vccd1 vccd1 _11603_/B sky130_fd_sc_hd__nor2_1
X_15370_ _15370_/A vssd1 vssd1 vccd1 vccd1 _15423_/C sky130_fd_sc_hd__clkbuf_1
X_12582_ _12582_/A _12582_/B vssd1 vssd1 vccd1 vccd1 _12589_/B sky130_fd_sc_hd__or2_1
XFILLER_106_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_208_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_196_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_184_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_180_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14321_ _14321_/A _14321_/B vssd1 vssd1 vccd1 vccd1 _14322_/B sky130_fd_sc_hd__or2_1
XFILLER_157_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11533_ _11522_/A _11532_/Y _12285_/C _11530_/A _19031_/Q vssd1 vssd1 vccd1 vccd1
+ _11534_/B sky130_fd_sc_hd__o2111a_1
XFILLER_184_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_1319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17040_ _17096_/A vssd1 vssd1 vccd1 vccd1 _17040_/X sky130_fd_sc_hd__clkbuf_2
X_11464_ _11478_/A _12340_/A _12340_/B _11828_/B vssd1 vssd1 vccd1 vccd1 _11464_/X
+ sky130_fd_sc_hd__a31o_1
X_14252_ _14257_/B _14252_/B vssd1 vssd1 vccd1 vccd1 _14305_/B sky130_fd_sc_hd__nor2_1
XFILLER_137_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13203_ _13203_/A vssd1 vssd1 vccd1 vccd1 _18057_/D sky130_fd_sc_hd__clkbuf_1
X_10415_ _10923_/S _10415_/B vssd1 vssd1 vccd1 vccd1 _10415_/Y sky130_fd_sc_hd__nand2_1
X_11395_ _11508_/C vssd1 vssd1 vccd1 vccd1 _11683_/A sky130_fd_sc_hd__clkbuf_2
X_14183_ _12027_/D _14120_/X _14152_/X _14167_/X _14182_/X vssd1 vssd1 vccd1 vccd1
+ _14183_/X sky130_fd_sc_hd__a2111o_4
XFILLER_109_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_1_1_wb_clk_i clkbuf_1_1_1_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_2_3_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_180_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10346_ _14260_/B _10343_/X _10345_/X _09916_/X vssd1 vssd1 vccd1 vccd1 _10346_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_124_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13134_ _13140_/A _18027_/Q vssd1 vssd1 vccd1 vccd1 _13135_/A sky130_fd_sc_hd__and2_1
XFILLER_140_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18991_ _18991_/CLK _18991_/D vssd1 vssd1 vccd1 vccd1 _18991_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_152_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_112_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13065_ _13394_/D _12776_/X _13064_/Y _13037_/X vssd1 vssd1 vccd1 vccd1 _17998_/D
+ sky130_fd_sc_hd__o211a_1
X_17942_ _18997_/CLK _17942_/D vssd1 vssd1 vccd1 vccd1 _17942_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_79_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_215_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10277_ _09198_/B _09193_/B _10286_/S vssd1 vssd1 vccd1 vccd1 _10277_/X sky130_fd_sc_hd__mux2_1
XFILLER_155_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12016_ _12025_/A _12016_/B vssd1 vssd1 vccd1 vccd1 _12016_/Y sky130_fd_sc_hd__nand2_1
XFILLER_79_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_215_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17873_ _19030_/CLK _17873_/D vssd1 vssd1 vccd1 vccd1 _17873_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_26_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_1366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16824_ _16866_/A _17425_/B _16866_/C vssd1 vssd1 vccd1 vccd1 _16824_/X sky130_fd_sc_hd__or3_1
XFILLER_207_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16755_ _16755_/A _16755_/B vssd1 vssd1 vccd1 vccd1 _16755_/Y sky130_fd_sc_hd__nand2_1
XFILLER_24_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_4_0_0_wb_clk_i clkbuf_4_1_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_5_1_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_2
X_13967_ _18442_/Q _13663_/X _13965_/X _13966_/X vssd1 vssd1 vccd1 vccd1 _13967_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_65_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15706_ _18542_/Q _18506_/Q _15714_/S vssd1 vssd1 vccd1 vccd1 _15706_/X sky130_fd_sc_hd__mux2_1
XFILLER_206_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12918_ _17969_/Q _12913_/X _12917_/Y vssd1 vssd1 vccd1 vccd1 _17969_/D sky130_fd_sc_hd__o21a_1
XFILLER_222_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16686_ _16699_/A _16686_/B vssd1 vssd1 vccd1 vccd1 _16686_/Y sky130_fd_sc_hd__nand2_1
X_13898_ _18532_/Q _13739_/X _13703_/A _18547_/Q vssd1 vssd1 vccd1 vccd1 _13898_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_179_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18425_ _18434_/CLK _18425_/D vssd1 vssd1 vccd1 vccd1 _18425_/Q sky130_fd_sc_hd__dfxtp_4
X_15637_ _18525_/Q _18489_/Q _15642_/S vssd1 vssd1 vccd1 vccd1 _15637_/X sky130_fd_sc_hd__mux2_1
XFILLER_206_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12849_ _12849_/A vssd1 vssd1 vccd1 vccd1 _17947_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_34_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_221_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18356_ _18356_/CLK _18356_/D vssd1 vssd1 vccd1 vccd1 _18356_/Q sky130_fd_sc_hd__dfxtp_2
X_15568_ _15568_/A vssd1 vssd1 vccd1 vccd1 _15586_/S sky130_fd_sc_hd__clkbuf_2
XTAP_1490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17307_ _18924_/Q _18888_/Q _17317_/S vssd1 vssd1 vccd1 vccd1 _17307_/X sky130_fd_sc_hd__mux2_1
XFILLER_119_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14519_ _18230_/Q _14515_/Y _14518_/X vssd1 vssd1 vccd1 vccd1 _18230_/D sky130_fd_sc_hd__o21ba_1
X_18287_ _18317_/CLK _18287_/D vssd1 vssd1 vccd1 vccd1 _18287_/Q sky130_fd_sc_hd__dfxtp_2
X_15499_ _18491_/Q _18455_/Q _15514_/S vssd1 vssd1 vccd1 vccd1 _15499_/X sky130_fd_sc_hd__mux2_1
XFILLER_175_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17238_ _17240_/B _17236_/X _17237_/Y _17219_/X vssd1 vssd1 vccd1 vccd1 _18871_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_70_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17169_ _17213_/A _17169_/B vssd1 vssd1 vccd1 vccd1 _17169_/Y sky130_fd_sc_hd__nand2_1
XFILLER_127_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_157_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_131_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09991_ _09991_/A vssd1 vssd1 vccd1 vccd1 _10103_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_157_1266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08942_ input1/X vssd1 vssd1 vccd1 vccd1 _08967_/A sky130_fd_sc_hd__buf_4
X_19096__67 vssd1 vssd1 vccd1 vccd1 _19096__67/HI _19204_/A sky130_fd_sc_hd__conb_1
XFILLER_88_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_229_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_225_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09425_ _09222_/Y _09454_/B _09425_/C vssd1 vssd1 vccd1 vccd1 _09482_/A sky130_fd_sc_hd__and3b_1
XFILLER_13_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_205_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09356_ _18278_/Q _18277_/Q _18276_/Q vssd1 vssd1 vccd1 vccd1 _09360_/A sky130_fd_sc_hd__or3_2
XFILLER_139_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_212_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_178_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_139_wb_clk_i clkbuf_5_27_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18350_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_205_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09287_ _09287_/A _09287_/B _09287_/C _09287_/D vssd1 vssd1 vccd1 vccd1 _09288_/C
+ sky130_fd_sc_hd__and4_1
XFILLER_201_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_1243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_1363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10200_ _10246_/A _10246_/B vssd1 vssd1 vccd1 vccd1 _10210_/A sky130_fd_sc_hd__xnor2_1
XFILLER_134_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11180_ _11181_/A _11184_/C vssd1 vssd1 vccd1 vccd1 _11185_/B sky130_fd_sc_hd__and2_1
XFILLER_107_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_1366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10131_ _10131_/A _10131_/B vssd1 vssd1 vccd1 vccd1 _10131_/Y sky130_fd_sc_hd__nor2_1
XFILLER_171_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_216_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10062_ _09181_/B _10009_/A _10061_/X vssd1 vssd1 vccd1 vccd1 _10065_/B sky130_fd_sc_hd__a21o_1
XTAP_5734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_173_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14870_ _14875_/B _14867_/X _14869_/X _14859_/X vssd1 vssd1 vccd1 vccd1 _18306_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_87_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13821_ _18576_/Q _13585_/A _13781_/X _18567_/Q _13820_/X vssd1 vssd1 vccd1 vccd1
+ _13821_/X sky130_fd_sc_hd__a221o_1
XFILLER_47_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_141_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16540_ _16538_/B _16537_/X _16538_/Y _16539_/X vssd1 vssd1 vccd1 vccd1 _18704_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_95_1334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13752_ _13752_/A vssd1 vssd1 vccd1 vccd1 _13752_/X sky130_fd_sc_hd__clkbuf_4
XINSDIODE2_108 _13954_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_216_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10964_ _10953_/X _10959_/X _10963_/X _09657_/X vssd1 vssd1 vccd1 vccd1 _10964_/X
+ sky130_fd_sc_hd__o31a_1
XINSDIODE2_119 _17471_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_231_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12703_ _12698_/Y _12702_/X _12522_/A vssd1 vssd1 vccd1 vccd1 _12707_/C sky130_fd_sc_hd__a21o_1
X_16471_ _16507_/A _16475_/B vssd1 vssd1 vccd1 vccd1 _16471_/Y sky130_fd_sc_hd__nand2_1
X_13683_ _18552_/Q _13573_/A _13676_/X _13682_/X vssd1 vssd1 vccd1 vccd1 _13683_/X
+ sky130_fd_sc_hd__a211o_2
XFILLER_16_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10895_ _10895_/A _10966_/B _10895_/C vssd1 vssd1 vccd1 vccd1 _10895_/X sky130_fd_sc_hd__and3_1
X_18210_ _18213_/CLK _18210_/D vssd1 vssd1 vccd1 vccd1 _18210_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_223_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15422_ _16935_/A vssd1 vssd1 vccd1 vccd1 _16021_/B sky130_fd_sc_hd__buf_2
XFILLER_188_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_203_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19190_ _19190_/A _08990_/Y vssd1 vssd1 vccd1 vccd1 io_out[28] sky130_fd_sc_hd__ebufn_8
X_12634_ _12627_/B _12569_/X _12632_/X _12633_/Y _12621_/X vssd1 vssd1 vccd1 vccd1
+ _17927_/D sky130_fd_sc_hd__a221o_1
XFILLER_169_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_223_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18141_ _18147_/CLK _18141_/D vssd1 vssd1 vccd1 vccd1 _18141_/Q sky130_fd_sc_hd__dfxtp_1
X_15353_ _15352_/B _15351_/X _15352_/Y _15340_/X vssd1 vssd1 vccd1 vccd1 _18422_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_129_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12565_ _12556_/A _12564_/X _12556_/B _12554_/B vssd1 vssd1 vccd1 vccd1 _12565_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_196_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14304_ _14275_/X _14298_/X _14303_/X _14270_/X vssd1 vssd1 vccd1 vccd1 _18176_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_102_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11516_ _11530_/B _11338_/A _11515_/Y vssd1 vssd1 vccd1 vccd1 _11516_/X sky130_fd_sc_hd__a21o_1
X_18072_ _18072_/CLK _18072_/D vssd1 vssd1 vccd1 vccd1 _18072_/Q sky130_fd_sc_hd__dfxtp_1
X_15284_ _15286_/B _15281_/X _15282_/Y _15283_/X vssd1 vssd1 vccd1 vccd1 _18409_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_89_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12496_ _14504_/B _12496_/B _12496_/C vssd1 vssd1 vccd1 vccd1 _12497_/A sky130_fd_sc_hd__and3_1
XFILLER_221_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17023_ _17035_/A _17023_/B vssd1 vssd1 vccd1 vccd1 _17023_/Y sky130_fd_sc_hd__nand2_1
XFILLER_8_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14235_ _14332_/S vssd1 vssd1 vccd1 vccd1 _14260_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_171_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11447_ _11447_/A vssd1 vssd1 vccd1 vccd1 _11788_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_7_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11378_ _11323_/B _11339_/C _11388_/A vssd1 vssd1 vccd1 vccd1 _11378_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_4_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14166_ _18986_/Q _14015_/X _14027_/X _18977_/Q _14165_/X vssd1 vssd1 vccd1 vccd1
+ _14166_/X sky130_fd_sc_hd__a221o_1
XFILLER_113_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_217_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13117_ _13117_/A vssd1 vssd1 vccd1 vccd1 _18018_/D sky130_fd_sc_hd__clkbuf_1
XTAP_504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10329_ _09282_/A _09287_/B _09287_/C _09282_/C _09969_/X _09935_/X vssd1 vssd1 vccd1
+ vccd1 _10329_/X sky130_fd_sc_hd__mux4_1
XFILLER_152_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14097_ _18650_/Q _13848_/X _13858_/A _18641_/Q vssd1 vssd1 vccd1 vccd1 _14097_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18974_ _18977_/CLK _18974_/D vssd1 vssd1 vccd1 vccd1 _18974_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13048_ _17995_/Q _12783_/A _13025_/A _13041_/Y _13368_/A vssd1 vssd1 vccd1 vccd1
+ _13049_/B sky130_fd_sc_hd__a32o_1
X_17925_ _18991_/CLK _17925_/D vssd1 vssd1 vccd1 vccd1 _17925_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_78_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17856_ _19034_/CLK _17856_/D vssd1 vssd1 vccd1 vccd1 _17856_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_15_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_227_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16807_ _16807_/A _16963_/C vssd1 vssd1 vccd1 vccd1 _16815_/B sky130_fd_sc_hd__nor2_1
XFILLER_26_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17787_ _17817_/CLK _17787_/D vssd1 vssd1 vccd1 vccd1 _17787_/Q sky130_fd_sc_hd__dfxtp_1
X_14999_ _15292_/A _15136_/C vssd1 vssd1 vccd1 vccd1 _15012_/B sky130_fd_sc_hd__nor2_1
XFILLER_19_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16738_ _18790_/Q _18754_/Q _16742_/S vssd1 vssd1 vccd1 vccd1 _16738_/X sky130_fd_sc_hd__mux2_1
XFILLER_207_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_222_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16669_ _18736_/Q _16670_/B _16668_/Y _16659_/X vssd1 vssd1 vccd1 vccd1 _18736_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_50_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_223_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09210_ _18698_/Q _18697_/Q _18696_/Q vssd1 vssd1 vccd1 vccd1 _09214_/A sky130_fd_sc_hd__or3_4
XFILLER_61_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18408_ _18408_/CLK _18408_/D vssd1 vssd1 vccd1 vccd1 _18408_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_210_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_148_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_232_wb_clk_i clkbuf_5_0_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17901_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_203_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09141_ _18722_/Q _18721_/Q _18720_/Q vssd1 vssd1 vccd1 vccd1 _09143_/C sky130_fd_sc_hd__or3_4
XFILLER_37_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18339_ _18343_/CLK _18339_/D vssd1 vssd1 vccd1 vccd1 _18339_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_72_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09072_ _09072_/A _09081_/B _17829_/Q vssd1 vssd1 vccd1 vccd1 _09073_/A sky130_fd_sc_hd__and3_1
XFILLER_136_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_118_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09974_ _09974_/A vssd1 vssd1 vccd1 vccd1 _10356_/A sky130_fd_sc_hd__buf_4
XFILLER_170_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_1260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_229_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_198_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_225_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_214_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_213_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09408_ _09408_/A _09408_/B _09408_/C _09408_/D vssd1 vssd1 vccd1 vccd1 _09419_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_41_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10680_ _10680_/A vssd1 vssd1 vccd1 vccd1 _12089_/A sky130_fd_sc_hd__buf_6
XFILLER_185_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09339_ _09339_/A _09443_/A vssd1 vssd1 vccd1 vccd1 _09421_/A sky130_fd_sc_hd__or2_4
XFILLER_194_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12350_ _12352_/B _12200_/X _12346_/A vssd1 vssd1 vccd1 vccd1 _12350_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_217_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11301_ _11301_/A _11899_/C vssd1 vssd1 vccd1 vccd1 _11501_/C sky130_fd_sc_hd__or2_1
XFILLER_153_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12281_ _12517_/A _12281_/B vssd1 vssd1 vccd1 vccd1 _12282_/A sky130_fd_sc_hd__and2_1
XFILLER_5_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14020_ _18857_/Q _13588_/X _13861_/X _18872_/Q vssd1 vssd1 vccd1 vccd1 _14020_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_5_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11232_ _11232_/A _11232_/B _11232_/C vssd1 vssd1 vccd1 vccd1 _11234_/A sky130_fd_sc_hd__and3_1
XFILLER_153_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11163_ _17822_/Q _17817_/Q _11245_/A _17823_/Q vssd1 vssd1 vccd1 vccd1 _11164_/D
+ sky130_fd_sc_hd__or4b_2
XFILLER_49_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_36_wb_clk_i clkbuf_5_5_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18875_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_1_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10114_ _18118_/Q _10114_/B vssd1 vssd1 vccd1 vccd1 _10122_/B sky130_fd_sc_hd__xnor2_4
X_15971_ _16003_/A _15971_/B vssd1 vssd1 vccd1 vccd1 _15971_/Y sky130_fd_sc_hd__nand2_1
XTAP_5520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11094_ _11895_/A vssd1 vssd1 vccd1 vccd1 _11113_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_49_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_1333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17710_ _17710_/A vssd1 vssd1 vccd1 vccd1 _18992_/D sky130_fd_sc_hd__clkbuf_1
XTAP_5553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14922_ _14980_/A vssd1 vssd1 vccd1 vccd1 _14922_/X sky130_fd_sc_hd__clkbuf_2
X_10045_ _10010_/A _10034_/X _10042_/X _10044_/X vssd1 vssd1 vccd1 vccd1 _10045_/X
+ sky130_fd_sc_hd__a211o_1
XTAP_5564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18690_ _18693_/CLK _18690_/D vssd1 vssd1 vccd1 vccd1 _18690_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_5575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17641_ _18183_/Q vssd1 vssd1 vccd1 vccd1 _17641_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_75_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14853_ _15292_/A _14989_/C vssd1 vssd1 vccd1 vccd1 _14861_/B sky130_fd_sc_hd__nor2_2
XFILLER_5_1260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13804_ _18369_/Q _13616_/A _13730_/A _18372_/Q _13803_/X vssd1 vssd1 vccd1 vccd1
+ _13804_/X sky130_fd_sc_hd__a221o_1
XFILLER_91_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17572_ _17571_/X _17560_/Y _17561_/X _17562_/Y _18956_/Q vssd1 vssd1 vccd1 vccd1
+ _17573_/B sky130_fd_sc_hd__a32o_1
XFILLER_217_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14784_ _18322_/Q _18286_/Q _14787_/S vssd1 vssd1 vccd1 vccd1 _14784_/X sky130_fd_sc_hd__mux2_1
XFILLER_44_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11996_ _11983_/A _11983_/B _11979_/A vssd1 vssd1 vccd1 vccd1 _12041_/C sky130_fd_sc_hd__a21o_2
XFILLER_189_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16523_ _18700_/Q _16525_/B _16522_/Y _16519_/X vssd1 vssd1 vccd1 vccd1 _18700_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_32_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_204_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13735_ _13735_/A vssd1 vssd1 vccd1 vccd1 _13735_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_32_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10947_ _09397_/B _10069_/A _10940_/X _09365_/D _10944_/S vssd1 vssd1 vccd1 vccd1
+ _10947_/X sky130_fd_sc_hd__a221o_1
XFILLER_45_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_189_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_182_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_108_1216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_220_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16454_ _18720_/Q _18684_/Q _16470_/S vssd1 vssd1 vccd1 vccd1 _16454_/X sky130_fd_sc_hd__mux2_1
XFILLER_108_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13666_ _13715_/A vssd1 vssd1 vccd1 vccd1 _13666_/X sky130_fd_sc_hd__buf_8
XFILLER_147_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10878_ _09397_/C _10644_/A _10877_/X _10693_/X vssd1 vssd1 vccd1 vccd1 _10878_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_182_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15405_ _15403_/B _15402_/X _15403_/Y _15404_/X vssd1 vssd1 vccd1 vccd1 _18434_/D
+ sky130_fd_sc_hd__o211a_1
XPHY_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19173_ _19173_/A _09021_/Y vssd1 vssd1 vccd1 vccd1 io_out[11] sky130_fd_sc_hd__ebufn_8
X_12617_ _12600_/A _12600_/B _12600_/C _12610_/B _12598_/B vssd1 vssd1 vccd1 vccd1
+ _12618_/B sky130_fd_sc_hd__a311oi_2
X_16385_ _16503_/A vssd1 vssd1 vccd1 vccd1 _16434_/A sky130_fd_sc_hd__dlymetal6s2s_1
XPHY_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13597_ _13706_/A vssd1 vssd1 vccd1 vccd1 _13630_/A sky130_fd_sc_hd__buf_8
XFILLER_157_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_223_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18124_ _18130_/CLK _18124_/D vssd1 vssd1 vccd1 vccd1 _18124_/Q sky130_fd_sc_hd__dfxtp_1
X_15336_ _15339_/B _15334_/X _15335_/Y _15315_/X vssd1 vssd1 vccd1 vccd1 _18418_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_185_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12548_ _12708_/A vssd1 vssd1 vccd1 vccd1 _12548_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_184_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_172_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18055_ _18068_/CLK _18055_/D vssd1 vssd1 vccd1 vccd1 _18055_/Q sky130_fd_sc_hd__dfxtp_1
X_15267_ _18441_/Q _18405_/Q _15267_/S vssd1 vssd1 vccd1 vccd1 _15267_/X sky130_fd_sc_hd__mux2_1
X_12479_ _12475_/Y _12476_/X _12499_/D _12484_/A _12472_/A vssd1 vssd1 vccd1 vccd1
+ _17907_/D sky130_fd_sc_hd__o311a_1
XFILLER_6_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17006_ _17032_/A _17010_/B vssd1 vssd1 vccd1 vccd1 _17006_/Y sky130_fd_sc_hd__nand2_1
X_14218_ _14295_/A vssd1 vssd1 vccd1 vccd1 _14335_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_193_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15198_ _18423_/Q _18387_/Q _15198_/S vssd1 vssd1 vccd1 vccd1 _15198_/X sky130_fd_sc_hd__mux2_1
XFILLER_125_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14149_ _18563_/Q _14017_/A _14145_/X _14148_/X vssd1 vssd1 vccd1 vccd1 _14149_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_119_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19066__37 vssd1 vssd1 vccd1 vccd1 _19066__37/HI _19160_/A sky130_fd_sc_hd__conb_1
X_18957_ _18959_/CLK _18957_/D vssd1 vssd1 vccd1 vccd1 _18957_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_67_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17908_ _19034_/CLK _17908_/D vssd1 vssd1 vccd1 vccd1 _17908_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_100_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09690_ _10600_/B _09676_/X _09677_/X _09678_/X _09683_/X _09689_/X vssd1 vssd1 vccd1
+ vccd1 _09691_/B sky130_fd_sc_hd__mux4_1
X_18888_ _18893_/CLK _18888_/D vssd1 vssd1 vccd1 vccd1 _18888_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_66_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17839_ _17890_/CLK _17839_/D vssd1 vssd1 vccd1 vccd1 _17839_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_55_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_215_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_228_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_1362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_207_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_1321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_212_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_222_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_223_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09124_ _18830_/Q _18829_/Q _18828_/Q vssd1 vssd1 vccd1 vccd1 _09126_/C sky130_fd_sc_hd__or3_4
XFILLER_182_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_148_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09055_ _09058_/A vssd1 vssd1 vccd1 vccd1 _09055_/Y sky130_fd_sc_hd__inv_2
XFILLER_198_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_194_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_1208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09957_ _10348_/A vssd1 vssd1 vccd1 vccd1 _09958_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_77_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09888_ _10370_/S _09979_/A vssd1 vssd1 vccd1 vccd1 _09889_/A sky130_fd_sc_hd__nor2_2
XTAP_890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_100_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19080__51 vssd1 vssd1 vccd1 vccd1 _19080__51/HI _19188_/A sky130_fd_sc_hd__conb_1
XFILLER_72_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11850_ _11850_/A _11850_/B _11850_/C _11850_/D vssd1 vssd1 vccd1 vccd1 _11850_/X
+ sky130_fd_sc_hd__or4_1
XTAP_2724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_154_wb_clk_i _18102_/CLK vssd1 vssd1 vccd1 vccd1 _18126_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_2746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10801_ _10799_/X _10800_/X _10801_/S vssd1 vssd1 vccd1 vccd1 _10801_/X sky130_fd_sc_hd__mux2_1
XFILLER_92_1304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11781_ _11781_/A _11781_/B vssd1 vssd1 vccd1 vccd1 _11781_/Y sky130_fd_sc_hd__nor2_1
XTAP_2779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_202_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13520_ _13741_/A vssd1 vssd1 vccd1 vccd1 _13594_/A sky130_fd_sc_hd__buf_2
XFILLER_159_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10732_ _12100_/A _12099_/A vssd1 vssd1 vccd1 vccd1 _10733_/A sky130_fd_sc_hd__and2b_2
XFILLER_207_1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_185_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13451_ _13452_/A _13452_/B _13447_/X _13450_/X vssd1 vssd1 vccd1 vccd1 _13451_/X
+ sky130_fd_sc_hd__a2bb2o_1
X_10663_ _10701_/A vssd1 vssd1 vccd1 vccd1 _10664_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_142_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_1260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_220_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12402_ _12409_/B _12403_/C _17897_/Q vssd1 vssd1 vccd1 vccd1 _12414_/A sky130_fd_sc_hd__o21a_1
XFILLER_40_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16170_ _18652_/Q _18616_/Q _16170_/S vssd1 vssd1 vccd1 vccd1 _16170_/X sky130_fd_sc_hd__mux2_1
XFILLER_185_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10594_ _09720_/A _10588_/X _10593_/X _10895_/A vssd1 vssd1 vccd1 vccd1 _10594_/X
+ sky130_fd_sc_hd__a22o_1
X_13382_ _09844_/A _11040_/X _11035_/B _13381_/X _13379_/B vssd1 vssd1 vccd1 vccd1
+ _18113_/D sky130_fd_sc_hd__o2111a_1
XFILLER_182_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_182_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15121_ _18405_/Q _18369_/Q _15121_/S vssd1 vssd1 vccd1 vccd1 _15121_/X sky130_fd_sc_hd__mux2_1
X_12333_ _17884_/Q _13066_/B _12333_/C vssd1 vssd1 vccd1 vccd1 _12334_/A sky130_fd_sc_hd__and3_1
XFILLER_5_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_177_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15052_ _18387_/Q _18351_/Q _15052_/S vssd1 vssd1 vccd1 vccd1 _15052_/X sky130_fd_sc_hd__mux2_1
XFILLER_126_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12264_ _12264_/A vssd1 vssd1 vccd1 vccd1 _17865_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_123_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14003_ _18940_/Q _13670_/X _13766_/A _18916_/Q vssd1 vssd1 vccd1 vccd1 _14003_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_107_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11215_ _17816_/Q _11215_/B vssd1 vssd1 vccd1 vccd1 _11224_/C sky130_fd_sc_hd__and2_1
X_12195_ _17911_/Q _17902_/Q _17901_/Q _17898_/Q vssd1 vssd1 vccd1 vccd1 _12197_/C
+ sky130_fd_sc_hd__or4_1
XFILLER_107_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18811_ _18811_/CLK _18811_/D vssd1 vssd1 vccd1 vccd1 _18811_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_6040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11146_ _11922_/A vssd1 vssd1 vccd1 vccd1 _11784_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_68_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_1272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15954_ _16000_/A _15960_/B vssd1 vssd1 vccd1 vccd1 _15954_/Y sky130_fd_sc_hd__nand2_1
X_18742_ _18743_/CLK _18742_/D vssd1 vssd1 vccd1 vccd1 _18742_/Q sky130_fd_sc_hd__dfxtp_2
X_11077_ _11368_/A _11232_/A _11091_/S vssd1 vssd1 vccd1 vccd1 _11078_/A sky130_fd_sc_hd__mux2_1
XTAP_5350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14905_ _18351_/Q _18315_/Q _14905_/S vssd1 vssd1 vccd1 vccd1 _14905_/X sky130_fd_sc_hd__mux2_1
XFILLER_37_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_1204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10028_ _10893_/S vssd1 vssd1 vccd1 vccd1 _10029_/S sky130_fd_sc_hd__clkbuf_4
X_18673_ _18677_/CLK _18673_/D vssd1 vssd1 vccd1 vccd1 _18673_/Q sky130_fd_sc_hd__dfxtp_4
XTAP_5394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15885_ _15885_/A vssd1 vssd1 vccd1 vccd1 _15938_/A sky130_fd_sc_hd__clkbuf_4
XTAP_4660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_224_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14836_ _14838_/B _14834_/X _14835_/Y _14819_/X vssd1 vssd1 vccd1 vccd1 _18298_/D
+ sky130_fd_sc_hd__o211a_1
X_17624_ _17623_/Y _17604_/X _17591_/X vssd1 vssd1 vccd1 vccd1 _17624_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_149_1338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17555_ _17548_/Y _17552_/X _18952_/Q vssd1 vssd1 vccd1 vccd1 _17555_/X sky130_fd_sc_hd__a21o_1
X_14767_ _14814_/A _14767_/B vssd1 vssd1 vccd1 vccd1 _14767_/Y sky130_fd_sc_hd__nand2_1
X_11979_ _11979_/A vssd1 vssd1 vccd1 vccd1 _12025_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_204_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16506_ _18733_/Q _18697_/Q _16509_/S vssd1 vssd1 vccd1 vccd1 _16506_/X sky130_fd_sc_hd__mux2_1
XFILLER_205_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13718_ _18246_/Q _13715_/X _13513_/A _18240_/Q _13717_/X vssd1 vssd1 vccd1 vccd1
+ _13718_/X sky130_fd_sc_hd__a221o_1
XFILLER_177_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17486_ _17509_/A _17489_/B vssd1 vssd1 vccd1 vccd1 _17486_/Y sky130_fd_sc_hd__nand2_1
XFILLER_220_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14698_ _15649_/A vssd1 vssd1 vccd1 vccd1 _14948_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_108_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_220_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16437_ _16456_/A vssd1 vssd1 vccd1 vccd1 _16437_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_19225_ _19225_/A _08931_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[25] sky130_fd_sc_hd__ebufn_8
XFILLER_20_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13649_ _13649_/A _13649_/B _13649_/C vssd1 vssd1 vccd1 vccd1 _13649_/X sky130_fd_sc_hd__and3_2
XFILLER_82_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_192_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19156_ _19156_/A _08951_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[26] sky130_fd_sc_hd__ebufn_8
X_16368_ _16807_/A _16504_/C vssd1 vssd1 vccd1 vccd1 _16378_/B sky130_fd_sc_hd__nor2_1
XFILLER_160_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18107_ _18130_/CLK _18107_/D vssd1 vssd1 vccd1 vccd1 _18107_/Q sky130_fd_sc_hd__dfxtp_2
X_15319_ _15578_/A vssd1 vssd1 vccd1 vccd1 _15373_/A sky130_fd_sc_hd__buf_2
XFILLER_9_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16299_ _16310_/A _16736_/B _16333_/C vssd1 vssd1 vccd1 vccd1 _16299_/X sky130_fd_sc_hd__or3_1
XFILLER_195_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_1339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18038_ _18094_/CLK _18038_/D vssd1 vssd1 vccd1 vccd1 _18038_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_195_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_126_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09811_ _12106_/A _12106_/B vssd1 vssd1 vccd1 vccd1 _10605_/A sky130_fd_sc_hd__nor2_2
XFILLER_98_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_140_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09742_ _09742_/A _09742_/B vssd1 vssd1 vccd1 vccd1 _09800_/A sky130_fd_sc_hd__xnor2_1
XFILLER_39_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09673_ _10041_/A vssd1 vssd1 vccd1 vccd1 _10962_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_39_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_223_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_4_13_0_wb_clk_i clkbuf_3_6_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_5_27_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_10_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_202_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09107_ _18755_/Q _18754_/Q _18753_/Q vssd1 vssd1 vccd1 vccd1 _09109_/C sky130_fd_sc_hd__or3_4
XFILLER_148_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09038_ _09040_/A vssd1 vssd1 vccd1 vccd1 _09038_/Y sky130_fd_sc_hd__inv_2
XFILLER_136_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11000_ _17823_/Q vssd1 vssd1 vccd1 vccd1 _11892_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_137_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12951_ _12951_/A _12951_/B vssd1 vssd1 vccd1 vccd1 _12951_/Y sky130_fd_sc_hd__nand2_1
XFILLER_46_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11902_ _12021_/A _11927_/A _11930_/B _17794_/Q vssd1 vssd1 vccd1 vccd1 _11947_/A
+ sky130_fd_sc_hd__a31o_1
XFILLER_73_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15670_ _15691_/A _15673_/B vssd1 vssd1 vccd1 vccd1 _15670_/Y sky130_fd_sc_hd__nand2_1
XFILLER_206_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12882_ _17957_/Q _12881_/B _12854_/X vssd1 vssd1 vccd1 vccd1 _12883_/B sky130_fd_sc_hd__o21ai_1
XTAP_3266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14621_ _18172_/Q _18171_/Q vssd1 vssd1 vccd1 vccd1 _14660_/B sky130_fd_sc_hd__or2b_1
XTAP_2543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11833_ _11393_/X _11374_/X _11828_/Y vssd1 vssd1 vccd1 vccd1 _11833_/X sky130_fd_sc_hd__o21a_1
XTAP_2554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17340_ _17376_/A _17483_/B _17376_/C vssd1 vssd1 vccd1 vccd1 _17340_/X sky130_fd_sc_hd__or3_1
X_14552_ _14690_/B _15156_/A vssd1 vssd1 vccd1 vccd1 _14559_/B sky130_fd_sc_hd__nor2_2
XFILLER_14_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11764_ _11764_/A _11770_/C vssd1 vssd1 vccd1 vccd1 _11764_/Y sky130_fd_sc_hd__nand2_1
XTAP_1864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13503_ _13677_/A vssd1 vssd1 vccd1 vccd1 _13719_/A sky130_fd_sc_hd__buf_6
XFILLER_18_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10715_ _09093_/A _09093_/B _09098_/C _09103_/B _10738_/A _10660_/X vssd1 vssd1 vccd1
+ vccd1 _10715_/X sky130_fd_sc_hd__mux4_2
XTAP_1897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17271_ _17318_/A _17415_/B _17318_/C vssd1 vssd1 vccd1 vccd1 _17271_/X sky130_fd_sc_hd__or3_1
XFILLER_186_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14483_ _18216_/Q _14491_/B vssd1 vssd1 vccd1 vccd1 _14484_/A sky130_fd_sc_hd__and2_1
X_11695_ _11689_/Y _11691_/Y _11709_/B _11694_/X _11689_/A vssd1 vssd1 vccd1 vccd1
+ _11696_/B sky130_fd_sc_hd__a32o_1
XFILLER_105_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19010_ _19029_/CLK _19010_/D vssd1 vssd1 vccd1 vccd1 _19010_/Q sky130_fd_sc_hd__dfxtp_1
X_16222_ _16807_/A _16358_/C vssd1 vssd1 vccd1 vccd1 _16229_/B sky130_fd_sc_hd__nor2_2
XFILLER_13_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13434_ _13434_/A _13434_/B _13434_/C vssd1 vssd1 vccd1 vccd1 _13436_/B sky130_fd_sc_hd__or3_1
XFILLER_179_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10646_ _10770_/A vssd1 vssd1 vccd1 vccd1 _10668_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_42_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16153_ _16909_/A vssd1 vssd1 vccd1 vccd1 _16749_/B sky130_fd_sc_hd__buf_4
X_13365_ _18106_/Q _13363_/Y _17704_/B _09509_/Y vssd1 vssd1 vccd1 vccd1 _18106_/D
+ sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_51_wb_clk_i clkbuf_5_5_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18860_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_10577_ _10090_/S _10574_/X _10576_/X _10041_/A vssd1 vssd1 vccd1 vccd1 _10577_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_10_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15104_ _15107_/B _15100_/X _15101_/Y _15103_/X vssd1 vssd1 vccd1 vccd1 _18364_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_170_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12316_ _17884_/Q _12316_/B _12316_/C vssd1 vssd1 vccd1 vccd1 _12316_/X sky130_fd_sc_hd__or3_1
XFILLER_5_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16084_ _16835_/A vssd1 vssd1 vccd1 vccd1 _16689_/A sky130_fd_sc_hd__buf_8
XFILLER_115_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13296_ _18069_/Q _18068_/Q _18071_/Q _18070_/Q vssd1 vssd1 vccd1 vccd1 _13297_/C
+ sky130_fd_sc_hd__or4_1
XFILLER_5_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15035_ _15038_/B _15033_/X _15034_/Y _15026_/X vssd1 vssd1 vccd1 vccd1 _18346_/D
+ sky130_fd_sc_hd__o211a_1
X_12247_ _11673_/A _11672_/B _12246_/Y _12258_/C _11639_/A vssd1 vssd1 vccd1 vccd1
+ _12248_/B sky130_fd_sc_hd__a32o_1
XFILLER_64_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_229_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12178_ _14436_/A vssd1 vssd1 vccd1 vccd1 _12178_/X sky130_fd_sc_hd__buf_4
XFILLER_3_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11129_ _11129_/A vssd1 vssd1 vccd1 vccd1 _17799_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_68_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_228_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16986_ _17012_/A vssd1 vssd1 vccd1 vccd1 _17109_/C sky130_fd_sc_hd__buf_2
XFILLER_111_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_209_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18725_ _18738_/CLK _18725_/D vssd1 vssd1 vccd1 vccd1 _18725_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_7_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_231_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15937_ _18598_/Q _18562_/Q _15937_/S vssd1 vssd1 vccd1 vccd1 _15937_/X sky130_fd_sc_hd__mux2_1
XTAP_5180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15868_ _18582_/Q _18546_/Q _15879_/S vssd1 vssd1 vccd1 vccd1 _15868_/X sky130_fd_sc_hd__mux2_1
X_18656_ _18658_/CLK _18656_/D vssd1 vssd1 vccd1 vccd1 _18656_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_4490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14819_ _14881_/A vssd1 vssd1 vccd1 vccd1 _14819_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_17607_ _17610_/A _17607_/B vssd1 vssd1 vccd1 vccd1 _17608_/A sky130_fd_sc_hd__and2_1
XFILLER_224_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15799_ _15799_/A _15946_/B _15811_/C vssd1 vssd1 vccd1 vccd1 _15799_/X sky130_fd_sc_hd__or3_1
X_18587_ _18590_/CLK _18587_/D vssd1 vssd1 vccd1 vccd1 _18587_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_196_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17538_ _17538_/A _17538_/B _17538_/C vssd1 vssd1 vccd1 vccd1 _17538_/X sky130_fd_sc_hd__or3_1
XFILLER_177_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_1335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_220_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17469_ _17512_/A _17469_/B vssd1 vssd1 vccd1 vccd1 _17469_/Y sky130_fd_sc_hd__nand2_1
XFILLER_123_1319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_225_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19208_ _19208_/A _08977_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[8] sky130_fd_sc_hd__ebufn_8
XFILLER_165_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19139_ _19139_/A _09037_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[9] sky130_fd_sc_hd__ebufn_8
XFILLER_195_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_218_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_218_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09725_ _09725_/A _09725_/B vssd1 vssd1 vccd1 vccd1 _09726_/B sky130_fd_sc_hd__xor2_2
XFILLER_68_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_216_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09656_ _12061_/A vssd1 vssd1 vccd1 vccd1 _09657_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_103_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19050__21 vssd1 vssd1 vccd1 vccd1 _19050__21/HI _19144_/A sky130_fd_sc_hd__conb_1
XFILLER_215_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_2_3_1_wb_clk_i clkbuf_2_3_1_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_7_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_216_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_215_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09587_ _09598_/S _09587_/B vssd1 vssd1 vccd1 vccd1 _09725_/B sky130_fd_sc_hd__xor2_2
XFILLER_203_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_184_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10500_ _09098_/C _09103_/B _09093_/A _09093_/B _10236_/A _10413_/X vssd1 vssd1 vccd1
+ vccd1 _10500_/X sky130_fd_sc_hd__mux4_2
XFILLER_128_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11480_ _11341_/A _12340_/A _11478_/Y _11489_/B vssd1 vssd1 vccd1 vccd1 _11480_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_7_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_184_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10431_ _09136_/D _09131_/D _09126_/C _09131_/B _10429_/X _10430_/X vssd1 vssd1 vccd1
+ vccd1 _10431_/X sky130_fd_sc_hd__mux4_1
Xclkbuf_5_2_0_wb_clk_i clkbuf_5_3_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _17864_/CLK
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_104_1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13150_ _13150_/A vssd1 vssd1 vccd1 vccd1 _18033_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_109_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10362_ _09098_/A _09093_/C _09103_/D _09098_/B _09937_/A _10349_/S vssd1 vssd1 vccd1
+ vccd1 _10362_/X sky130_fd_sc_hd__mux4_1
XFILLER_128_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12101_ _12101_/A _12101_/B vssd1 vssd1 vccd1 vccd1 _12103_/C sky130_fd_sc_hd__xnor2_1
X_10293_ _10293_/A _10600_/A vssd1 vssd1 vccd1 vccd1 _10293_/X sky130_fd_sc_hd__or2_1
XFILLER_124_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13081_ _13081_/A vssd1 vssd1 vccd1 vccd1 _18003_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_151_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12032_ _12032_/A _12089_/B vssd1 vssd1 vccd1 vccd1 _12032_/X sky130_fd_sc_hd__xor2_1
XFILLER_215_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_215_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16840_ _16866_/A _17437_/B _16866_/C vssd1 vssd1 vccd1 vccd1 _16840_/X sky130_fd_sc_hd__or3_1
XFILLER_77_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16771_ _16771_/A _16794_/B vssd1 vssd1 vccd1 vccd1 _16779_/B sky130_fd_sc_hd__nor2_2
XFILLER_24_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_1310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13983_ _18346_/Q _13749_/A _13979_/X _13982_/X vssd1 vssd1 vccd1 vccd1 _13983_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_150_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18510_ _18511_/CLK _18510_/D vssd1 vssd1 vccd1 vccd1 _18510_/Q sky130_fd_sc_hd__dfxtp_2
X_15722_ _16019_/A _15745_/B vssd1 vssd1 vccd1 vccd1 _15730_/B sky130_fd_sc_hd__nor2_1
XFILLER_24_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12934_ _11044_/B _12933_/A _12933_/Y _12318_/X vssd1 vssd1 vccd1 vccd1 _17970_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_3030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_1278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15653_ _15944_/A _15696_/B vssd1 vssd1 vccd1 vccd1 _15661_/B sky130_fd_sc_hd__nor2_2
X_18441_ _18473_/CLK _18441_/D vssd1 vssd1 vccd1 vccd1 _18441_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_2_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12865_ _17951_/Q _17952_/Q _12865_/C vssd1 vssd1 vccd1 vccd1 _12868_/B sky130_fd_sc_hd__and3_1
XFILLER_73_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14604_ _14604_/A _14606_/B vssd1 vssd1 vccd1 vccd1 _14604_/Y sky130_fd_sc_hd__nand2_1
XFILLER_2_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18372_ _18374_/CLK _18372_/D vssd1 vssd1 vccd1 vccd1 _18372_/Q sky130_fd_sc_hd__dfxtp_2
X_11816_ _17517_/A vssd1 vssd1 vccd1 vccd1 _11816_/X sky130_fd_sc_hd__buf_4
XTAP_2384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15584_ _15583_/B _15581_/X _15583_/Y _15575_/X vssd1 vssd1 vccd1 vccd1 _18476_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_1650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12796_ _17964_/Q vssd1 vssd1 vccd1 vccd1 _12796_/Y sky130_fd_sc_hd__inv_2
XTAP_2395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17323_ _17323_/A vssd1 vssd1 vccd1 vccd1 _17400_/A sky130_fd_sc_hd__buf_2
XFILLER_187_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14535_ _18183_/Q vssd1 vssd1 vccd1 vccd1 _15951_/A sky130_fd_sc_hd__inv_2
X_11747_ _11747_/A _11761_/B vssd1 vssd1 vccd1 vccd1 _11749_/B sky130_fd_sc_hd__xor2_2
XTAP_1694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_222_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17254_ _17536_/A _17254_/B vssd1 vssd1 vccd1 vccd1 _17263_/B sky130_fd_sc_hd__nor2_2
X_14466_ _14470_/C _14466_/B vssd1 vssd1 vccd1 vccd1 _18208_/D sky130_fd_sc_hd__nor2_1
X_11678_ _11374_/A _13429_/A _11635_/A _11257_/B _11652_/B vssd1 vssd1 vccd1 vccd1
+ _11845_/A sky130_fd_sc_hd__a2111o_2
X_16205_ _16794_/A _16205_/B vssd1 vssd1 vccd1 vccd1 _16217_/B sky130_fd_sc_hd__nor2_1
XFILLER_122_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13417_ _14507_/A _13417_/B vssd1 vssd1 vccd1 vccd1 _13418_/D sky130_fd_sc_hd__nand2_1
XFILLER_190_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17185_ _17193_/A _17473_/B _17234_/C vssd1 vssd1 vccd1 vccd1 _17185_/X sky130_fd_sc_hd__or3_1
X_10629_ _10629_/A vssd1 vssd1 vccd1 vccd1 _12958_/A sky130_fd_sc_hd__clkbuf_4
X_14397_ _17591_/A vssd1 vssd1 vccd1 vccd1 _14414_/A sky130_fd_sc_hd__buf_2
XFILLER_155_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16136_ _18645_/Q _18609_/Q _16145_/S vssd1 vssd1 vccd1 vccd1 _16136_/X sky130_fd_sc_hd__mux2_1
XFILLER_155_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13348_ _13348_/A _13389_/B vssd1 vssd1 vccd1 vccd1 _13348_/Y sky130_fd_sc_hd__nand2_1
XFILLER_170_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_192_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16067_ _16672_/A _16208_/C vssd1 vssd1 vccd1 vccd1 _16082_/B sky130_fd_sc_hd__nor2_2
XFILLER_5_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13279_ _19006_/Q _19005_/Q _19008_/Q _19007_/Q vssd1 vssd1 vccd1 vccd1 _13281_/A
+ sky130_fd_sc_hd__or4_1
XFILLER_45_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15018_ _18378_/Q _18342_/Q _15033_/S vssd1 vssd1 vccd1 vccd1 _15018_/X sky130_fd_sc_hd__mux2_1
XFILLER_102_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_229_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16969_ _16972_/B _16966_/X _16968_/Y _16964_/X vssd1 vssd1 vccd1 vccd1 _18805_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_110_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_231_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09510_ input2/X vssd1 vssd1 vccd1 vccd1 _12217_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_65_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18708_ _18708_/CLK _18708_/D vssd1 vssd1 vccd1 vccd1 _18708_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_224_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09441_ _09420_/A _09419_/Y _09450_/A vssd1 vssd1 vccd1 vccd1 _09441_/X sky130_fd_sc_hd__o21ba_1
X_18639_ _18641_/CLK _18639_/D vssd1 vssd1 vccd1 vccd1 _18639_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_25_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_224_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_220_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09372_ _18407_/Q _18406_/Q _18405_/Q vssd1 vssd1 vccd1 vccd1 _09376_/A sky130_fd_sc_hd__or3_4
XFILLER_36_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_220_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_220_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINSDIODE2_2 _08960_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_5916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_181_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_229_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_229_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_229_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09708_ _09708_/A vssd1 vssd1 vccd1 vccd1 _09709_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_216_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10980_ _12361_/A vssd1 vssd1 vccd1 vccd1 _15840_/A sky130_fd_sc_hd__buf_12
XFILLER_55_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09639_ _09669_/B _09639_/B vssd1 vssd1 vccd1 vccd1 _09640_/B sky130_fd_sc_hd__xnor2_4
XFILLER_55_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_188_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12650_ _12649_/A _12649_/B _12591_/X vssd1 vssd1 vccd1 vccd1 _12650_/X sky130_fd_sc_hd__o21a_1
XFILLER_169_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_231_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_208_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11601_ _17857_/Q _17856_/Q vssd1 vssd1 vccd1 vccd1 _11602_/B sky130_fd_sc_hd__or2_1
XFILLER_208_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12581_ _12561_/Y _12573_/A _12571_/X _12575_/B vssd1 vssd1 vccd1 vccd1 _12582_/B
+ sky130_fd_sc_hd__a31oi_4
XFILLER_23_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14320_ _14321_/A _14321_/B vssd1 vssd1 vccd1 vccd1 _14334_/A sky130_fd_sc_hd__nand2_1
XFILLER_12_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11532_ _12285_/B vssd1 vssd1 vccd1 vccd1 _11532_/Y sky130_fd_sc_hd__inv_2
XFILLER_157_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14251_ _14464_/A _14323_/C vssd1 vssd1 vccd1 vccd1 _14252_/B sky130_fd_sc_hd__nor2_1
X_11463_ _11479_/B _11463_/B vssd1 vssd1 vccd1 vccd1 _12340_/B sky130_fd_sc_hd__nand2_1
XFILLER_137_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13202_ _13208_/A _18058_/Q vssd1 vssd1 vccd1 vccd1 _13203_/A sky130_fd_sc_hd__and2_1
XFILLER_137_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10414_ _09209_/A _09219_/B _09214_/D _09214_/B _10496_/A _10413_/X vssd1 vssd1 vccd1
+ vccd1 _10415_/B sky130_fd_sc_hd__mux4_2
X_14182_ _13693_/Y _14174_/X _14181_/X _12042_/B _13416_/A vssd1 vssd1 vccd1 vccd1
+ _14182_/X sky130_fd_sc_hd__a221o_4
XFILLER_99_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11394_ _11374_/X _11384_/Y _11391_/Y _11393_/X vssd1 vssd1 vccd1 vccd1 _11394_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_136_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13133_ _13133_/A vssd1 vssd1 vccd1 vccd1 _18025_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_178_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10345_ _10356_/A _10345_/B vssd1 vssd1 vccd1 vccd1 _10345_/X sky130_fd_sc_hd__or2_1
XFILLER_139_1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18990_ _18991_/CLK _18990_/D vssd1 vssd1 vccd1 vccd1 _18990_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_79_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_124_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17941_ _18993_/CLK _17941_/D vssd1 vssd1 vccd1 vccd1 _17941_/Q sky130_fd_sc_hd__dfxtp_2
X_13064_ _13052_/X _13063_/Y _12786_/B vssd1 vssd1 vccd1 vccd1 _13064_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_152_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10276_ _10375_/S vssd1 vssd1 vccd1 vccd1 _10286_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_152_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_215_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_1334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12015_ _12015_/A _12015_/B vssd1 vssd1 vccd1 vccd1 _12015_/Y sky130_fd_sc_hd__nand2_1
X_17872_ _19030_/CLK _17872_/D vssd1 vssd1 vccd1 vccd1 _17872_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_79_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_215_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_215_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16823_ _16823_/A vssd1 vssd1 vccd1 vccd1 _17425_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_120_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_226_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13966_ _18430_/Q _13785_/X _13766_/X _18412_/Q vssd1 vssd1 vccd1 vccd1 _13966_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_171_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16754_ _18794_/Q _18758_/Q _16762_/S vssd1 vssd1 vccd1 vccd1 _16754_/X sky130_fd_sc_hd__mux2_1
XFILLER_150_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_206_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15705_ _15708_/B _15702_/X _15704_/Y _15700_/X vssd1 vssd1 vccd1 vccd1 _18505_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_62_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12917_ _17969_/Q _12913_/X _12888_/B vssd1 vssd1 vccd1 vccd1 _12917_/Y sky130_fd_sc_hd__a21boi_1
X_16685_ _18776_/Q _18740_/Q _16694_/S vssd1 vssd1 vccd1 vccd1 _16685_/X sky130_fd_sc_hd__mux2_1
X_13897_ _18625_/Q _13573_/A _13531_/A _18616_/Q _13896_/X vssd1 vssd1 vccd1 vccd1
+ _13897_/X sky130_fd_sc_hd__a221o_1
XFILLER_62_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18424_ _18434_/CLK _18424_/D vssd1 vssd1 vccd1 vccd1 _18424_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_61_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15636_ _15931_/A _15696_/B vssd1 vssd1 vccd1 vccd1 _15651_/B sky130_fd_sc_hd__nor2_2
XFILLER_221_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12848_ _12851_/B _12848_/B _12915_/B vssd1 vssd1 vccd1 vccd1 _12849_/A sky130_fd_sc_hd__and3b_1
XTAP_2170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_146_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15567_ _15570_/B _15565_/X _15566_/Y _15555_/X vssd1 vssd1 vccd1 vccd1 _18472_/D
+ sky130_fd_sc_hd__o211a_1
X_18355_ _18356_/CLK _18355_/D vssd1 vssd1 vccd1 vccd1 _18355_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_226_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12779_ _18003_/Q vssd1 vssd1 vccd1 vccd1 _13082_/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_1491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_203_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14518_ _18230_/Q _14515_/Y _14377_/A vssd1 vssd1 vccd1 vccd1 _14518_/X sky130_fd_sc_hd__a21o_1
X_17306_ _17446_/A _17351_/B vssd1 vssd1 vccd1 vccd1 _17314_/B sky130_fd_sc_hd__nor2_1
X_15498_ _15568_/A vssd1 vssd1 vccd1 vccd1 _15514_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_148_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18286_ _18317_/CLK _18286_/D vssd1 vssd1 vccd1 vccd1 _18286_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_31_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14449_ _14449_/A vssd1 vssd1 vccd1 vccd1 _18202_/D sky130_fd_sc_hd__clkbuf_1
X_17237_ _17273_/A _17240_/B vssd1 vssd1 vccd1 vccd1 _17237_/Y sky130_fd_sc_hd__nand2_1
XFILLER_163_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17168_ _17168_/A vssd1 vssd1 vccd1 vccd1 _17213_/A sky130_fd_sc_hd__buf_2
XFILLER_157_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16119_ _16130_/A _16123_/B vssd1 vssd1 vccd1 vccd1 _16119_/Y sky130_fd_sc_hd__nand2_1
XFILLER_6_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17099_ _18874_/Q _18838_/Q _17114_/S vssd1 vssd1 vccd1 vccd1 _17099_/X sky130_fd_sc_hd__mux2_1
X_09990_ _10102_/S vssd1 vssd1 vccd1 vccd1 _10003_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_89_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08941_ _08941_/A vssd1 vssd1 vccd1 vccd1 _08941_/Y sky130_fd_sc_hd__inv_2
XFILLER_103_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_229_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_231_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_225_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_231_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09424_ _09421_/A _09427_/A _09450_/B vssd1 vssd1 vccd1 vccd1 _09425_/C sky130_fd_sc_hd__o21ai_4
XFILLER_225_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_197_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09355_ _09355_/A _09355_/B _09355_/C vssd1 vssd1 vccd1 vccd1 _09427_/A sky130_fd_sc_hd__nand3_4
XFILLER_205_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_221_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_205_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09286_ _18848_/Q _18847_/Q _18846_/Q vssd1 vssd1 vccd1 vccd1 _09287_/D sky130_fd_sc_hd__or3_4
XFILLER_60_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_179_wb_clk_i clkbuf_5_10_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18035_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_119_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_118_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_108_wb_clk_i clkbuf_5_29_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18563_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_10_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10130_ _10440_/A _10440_/B vssd1 vssd1 vccd1 vccd1 _10441_/A sky130_fd_sc_hd__nor2_4
XFILLER_133_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10061_ _09165_/C _10040_/A _09999_/A _09198_/B _10060_/X vssd1 vssd1 vccd1 vccd1
+ _10061_/X sky130_fd_sc_hd__a221o_1
XFILLER_0_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_197_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_85_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13820_ _18570_/Q _13715_/A _13623_/A _18564_/Q vssd1 vssd1 vccd1 vccd1 _13820_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_169_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_229_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13751_ _18792_/Q _13560_/A _13715_/X _18786_/Q _13750_/X vssd1 vssd1 vccd1 vccd1
+ _13751_/X sky130_fd_sc_hd__a221o_1
XINSDIODE2_109 _14027_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10963_ _09711_/A _10960_/X _10962_/X _10940_/X vssd1 vssd1 vccd1 vccd1 _10963_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_21_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12702_ _12688_/A _12688_/B _12693_/A _12701_/X vssd1 vssd1 vccd1 vccd1 _12702_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_203_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16470_ _18724_/Q _18688_/Q _16470_/S vssd1 vssd1 vccd1 vccd1 _16470_/X sky130_fd_sc_hd__mux2_1
X_13682_ _18537_/Q _13596_/A _13586_/A _18540_/Q _13681_/X vssd1 vssd1 vccd1 vccd1
+ _13682_/X sky130_fd_sc_hd__a221o_1
XFILLER_231_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10894_ _09720_/A _10890_/X _10893_/X _12061_/A vssd1 vssd1 vccd1 vccd1 _10895_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_71_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15421_ _18474_/Q _18438_/Q _15435_/S vssd1 vssd1 vccd1 vccd1 _15421_/X sky130_fd_sc_hd__mux2_1
X_12633_ _12632_/A _12632_/B _12569_/A vssd1 vssd1 vccd1 vccd1 _12633_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_71_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_231_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_223_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15352_ _15375_/A _15352_/B vssd1 vssd1 vccd1 vccd1 _15352_/Y sky130_fd_sc_hd__nand2_1
XFILLER_169_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18140_ _18140_/CLK _18140_/D vssd1 vssd1 vccd1 vccd1 _18140_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_12_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_223_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12564_ _12564_/A _17919_/Q vssd1 vssd1 vccd1 vccd1 _12564_/X sky130_fd_sc_hd__or2_1
X_14303_ _14299_/X _14282_/X _14283_/X _14300_/X _15145_/A vssd1 vssd1 vccd1 vccd1
+ _14303_/X sky130_fd_sc_hd__a311o_1
XFILLER_141_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18071_ _18072_/CLK _18071_/D vssd1 vssd1 vccd1 vccd1 _18071_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_11_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11515_ _17872_/Q _12279_/A vssd1 vssd1 vccd1 vccd1 _11515_/Y sky130_fd_sc_hd__nor2_1
X_15283_ _15283_/A vssd1 vssd1 vccd1 vccd1 _15283_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_32_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12495_ _12495_/A _12495_/B _12495_/C _12495_/D vssd1 vssd1 vccd1 vccd1 _12496_/C
+ sky130_fd_sc_hd__nand4_1
X_17022_ _18854_/Q _18818_/Q _17026_/S vssd1 vssd1 vccd1 vccd1 _17022_/X sky130_fd_sc_hd__mux2_1
XFILLER_116_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14234_ _14323_/C _14463_/B vssd1 vssd1 vccd1 vccd1 _14234_/Y sky130_fd_sc_hd__nand2_1
XFILLER_221_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11446_ _11683_/A _11730_/B _11413_/Y _11429_/Y _11445_/X vssd1 vssd1 vccd1 vccd1
+ _11446_/X sky130_fd_sc_hd__a41o_1
XFILLER_137_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14165_ _18959_/Q _14017_/X _14161_/X _14164_/X vssd1 vssd1 vccd1 vccd1 _14165_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_217_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11377_ _11377_/A vssd1 vssd1 vccd1 vccd1 _11828_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_153_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13116_ _13118_/A _18019_/Q vssd1 vssd1 vccd1 vccd1 _13117_/A sky130_fd_sc_hd__and2_1
XFILLER_113_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10328_ _10320_/X _10327_/X _09981_/X vssd1 vssd1 vccd1 vccd1 _10328_/X sky130_fd_sc_hd__o21a_1
X_14096_ _18413_/Q _13539_/X _14090_/X _14095_/X vssd1 vssd1 vccd1 vccd1 _14096_/X
+ sky130_fd_sc_hd__a211o_1
XTAP_516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18973_ _18977_/CLK _18973_/D vssd1 vssd1 vccd1 vccd1 _18973_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_113_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13047_ _13047_/A vssd1 vssd1 vccd1 vccd1 _17994_/D sky130_fd_sc_hd__clkbuf_1
X_17924_ _18988_/CLK _17924_/D vssd1 vssd1 vccd1 vccd1 _17924_/Q sky130_fd_sc_hd__dfxtp_1
X_10259_ _10215_/A _10192_/B _10258_/X vssd1 vssd1 vccd1 vccd1 _11916_/B sky130_fd_sc_hd__o21ba_1
XFILLER_230_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17855_ _17891_/CLK _17855_/D vssd1 vssd1 vccd1 vccd1 _17855_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16806_ _16879_/A vssd1 vssd1 vccd1 vccd1 _16963_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_93_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17786_ _17817_/CLK _17786_/D vssd1 vssd1 vccd1 vccd1 _17786_/Q sky130_fd_sc_hd__dfxtp_1
X_14998_ _15064_/A vssd1 vssd1 vccd1 vccd1 _15136_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_47_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16737_ _16743_/B _16735_/X _16736_/X _16724_/X vssd1 vssd1 vccd1 vccd1 _18753_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_53_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13949_ _18505_/Q _13848_/A _13654_/X _18496_/Q _13948_/X vssd1 vssd1 vccd1 vccd1
+ _13949_/X sky130_fd_sc_hd__a221o_1
XFILLER_208_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_207_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16668_ _16695_/A _16670_/B vssd1 vssd1 vccd1 vccd1 _16668_/Y sky130_fd_sc_hd__nand2_1
XFILLER_201_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_210_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18407_ _18432_/CLK _18407_/D vssd1 vssd1 vccd1 vccd1 _18407_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_62_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15619_ _18485_/Q _15618_/B _15618_/Y _15616_/X vssd1 vssd1 vccd1 vccd1 _18485_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_210_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16599_ _16634_/A _16599_/B vssd1 vssd1 vccd1 vccd1 _16599_/Y sky130_fd_sc_hd__nand2_1
XFILLER_50_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09140_ _18707_/Q _18706_/Q _18705_/Q vssd1 vssd1 vccd1 vccd1 _09143_/B sky130_fd_sc_hd__or3_4
XFILLER_163_1271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18338_ _18373_/CLK _18338_/D vssd1 vssd1 vccd1 vccd1 _18338_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_37_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_6_wb_clk_i _17929_/CLK vssd1 vssd1 vccd1 vccd1 _18204_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_148_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09071_ _17837_/Q vssd1 vssd1 vccd1 vccd1 _09081_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_148_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18269_ _18275_/CLK _18269_/D vssd1 vssd1 vccd1 vccd1 _18269_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_190_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_201_wb_clk_i _18176_/CLK vssd1 vssd1 vccd1 vccd1 _18967_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_116_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_226_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_143_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09973_ _09381_/C _09945_/X _09972_/X _09923_/X vssd1 vssd1 vccd1 vccd1 _09973_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_131_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_226_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_217_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_225_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_214_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09407_ _18338_/Q _18337_/Q _18336_/Q vssd1 vssd1 vccd1 vccd1 _09408_/D sky130_fd_sc_hd__or3_1
XFILLER_38_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_1330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09338_ _09338_/A _09338_/B _09338_/C vssd1 vssd1 vccd1 vccd1 _09443_/A sky130_fd_sc_hd__and3_1
XFILLER_139_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_205_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09269_ _18986_/Q _18985_/Q _18984_/Q vssd1 vssd1 vccd1 vccd1 _09270_/D sky130_fd_sc_hd__or3_2
XFILLER_139_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11300_ _17793_/Q _17792_/Q _17794_/Q vssd1 vssd1 vccd1 vccd1 _11899_/C sky130_fd_sc_hd__or3b_4
XFILLER_193_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12280_ _12279_/Y _12279_/A _12289_/A vssd1 vssd1 vccd1 vccd1 _12281_/B sky130_fd_sc_hd__mux2_1
XFILLER_112_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11231_ _11231_/A _11231_/B vssd1 vssd1 vccd1 vccd1 _17819_/D sky130_fd_sc_hd__nor2_1
XFILLER_101_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11162_ _17824_/Q vssd1 vssd1 vccd1 vccd1 _11245_/A sky130_fd_sc_hd__inv_2
XFILLER_45_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10113_ _10113_/A vssd1 vssd1 vccd1 vccd1 _10122_/A sky130_fd_sc_hd__inv_2
XFILLER_110_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15970_ _18605_/Q _18569_/Q _15990_/S vssd1 vssd1 vccd1 vccd1 _15970_/X sky130_fd_sc_hd__mux2_1
XTAP_5510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11093_ _17793_/Q vssd1 vssd1 vccd1 vccd1 _12041_/A sky130_fd_sc_hd__buf_2
XFILLER_110_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_216_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14921_ _14932_/A _14924_/B vssd1 vssd1 vccd1 vccd1 _14921_/Y sky130_fd_sc_hd__nand2_1
X_10044_ _10044_/A _10044_/B vssd1 vssd1 vccd1 vccd1 _10044_/X sky130_fd_sc_hd__and2_1
XTAP_5554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_76_wb_clk_i clkbuf_5_21_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18641_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_5565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17640_ _17640_/A vssd1 vssd1 vccd1 vccd1 _17659_/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_5598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14852_ _14918_/A vssd1 vssd1 vccd1 vccd1 _14989_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_91_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_224_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_1272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13803_ _18345_/Q _13749_/A _13799_/X _13802_/X vssd1 vssd1 vccd1 vccd1 _13803_/X
+ sky130_fd_sc_hd__a211o_1
X_14783_ _14788_/B _14781_/X _14782_/X _14778_/X vssd1 vssd1 vccd1 vccd1 _18285_/D
+ sky130_fd_sc_hd__o211a_1
X_17571_ _18184_/Q vssd1 vssd1 vccd1 vccd1 _17571_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_63_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11995_ _13518_/B vssd1 vssd1 vccd1 vccd1 _12092_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_91_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16522_ _16572_/A _16525_/B vssd1 vssd1 vccd1 vccd1 _16522_/Y sky130_fd_sc_hd__nand2_1
X_13734_ _13734_/A vssd1 vssd1 vccd1 vccd1 _13734_/X sky130_fd_sc_hd__buf_4
XFILLER_182_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10946_ _09397_/D _10069_/X _10940_/X _09365_/B _10948_/S vssd1 vssd1 vccd1 vccd1
+ _10946_/X sky130_fd_sc_hd__a221o_1
XFILLER_56_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_205_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_1293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16453_ _16473_/A vssd1 vssd1 vccd1 vccd1 _16470_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_189_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13665_ _18873_/Q _13663_/X _13664_/X _18849_/Q vssd1 vssd1 vccd1 vccd1 _13665_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_220_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_182_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10877_ _10877_/A _10877_/B vssd1 vssd1 vccd1 vccd1 _10877_/X sky130_fd_sc_hd__or2_1
XFILLER_108_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_223_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_1299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15404_ _15404_/A vssd1 vssd1 vccd1 vccd1 _15404_/X sky130_fd_sc_hd__clkbuf_2
XPHY_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12616_ _12616_/A vssd1 vssd1 vccd1 vccd1 _12619_/A sky130_fd_sc_hd__inv_2
X_16384_ _18702_/Q _18666_/Q _16400_/S vssd1 vssd1 vccd1 vccd1 _16384_/X sky130_fd_sc_hd__mux2_1
X_19172_ _19172_/A _09020_/Y vssd1 vssd1 vccd1 vccd1 io_out[10] sky130_fd_sc_hd__ebufn_8
XPHY_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13596_ _13596_/A vssd1 vssd1 vccd1 vccd1 _13596_/X sky130_fd_sc_hd__clkbuf_4
XPHY_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15335_ _15373_/A _15339_/B vssd1 vssd1 vccd1 vccd1 _15335_/Y sky130_fd_sc_hd__nand2_1
XFILLER_8_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18123_ _18130_/CLK _18123_/D vssd1 vssd1 vccd1 vccd1 _18123_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_157_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12547_ _12544_/X _12556_/A _12542_/Y _12569_/A vssd1 vssd1 vccd1 vccd1 _12547_/Y
+ sky130_fd_sc_hd__a31oi_1
XFILLER_61_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15266_ _15266_/A _15277_/B vssd1 vssd1 vccd1 vccd1 _15275_/B sky130_fd_sc_hd__nor2_2
XFILLER_157_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18054_ _18068_/CLK _18054_/D vssd1 vssd1 vccd1 vccd1 _18054_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_144_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12478_ _12476_/X _12499_/D _12475_/Y vssd1 vssd1 vccd1 vccd1 _12484_/A sky130_fd_sc_hd__o21ai_1
X_17005_ _18850_/Q _18814_/Q _17005_/S vssd1 vssd1 vccd1 vccd1 _17005_/X sky130_fd_sc_hd__mux2_1
X_14217_ _18211_/Q _14196_/C _14211_/X _14342_/B _14342_/A vssd1 vssd1 vccd1 vccd1
+ _14295_/A sky130_fd_sc_hd__o311a_1
XFILLER_172_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11429_ _11415_/Y _11425_/Y _11428_/Y vssd1 vssd1 vccd1 vccd1 _11429_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_6_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15197_ _15197_/A _15229_/B vssd1 vssd1 vccd1 vccd1 _15206_/B sky130_fd_sc_hd__nor2_2
XFILLER_126_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14148_ _18587_/Q _13617_/A _14146_/X _14147_/X vssd1 vssd1 vccd1 vccd1 _14148_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_141_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14079_ _18707_/Q _13619_/X _14075_/X _14078_/X vssd1 vssd1 vccd1 vccd1 _14079_/X
+ sky130_fd_sc_hd__a211o_1
X_18956_ _18959_/CLK _18956_/D vssd1 vssd1 vccd1 vccd1 _18956_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_141_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17907_ _17907_/CLK _17907_/D vssd1 vssd1 vccd1 vccd1 _17907_/Q sky130_fd_sc_hd__dfxtp_1
X_18887_ _18893_/CLK _18887_/D vssd1 vssd1 vccd1 vccd1 _18887_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_230_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17838_ _17851_/CLK _17838_/D vssd1 vssd1 vccd1 vccd1 _17838_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_54_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_227_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_212_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_208_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17769_ _17769_/A vssd1 vssd1 vccd1 vccd1 _19027_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_78_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_228_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_1366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_223_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_206_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09123_ _18815_/Q _18814_/Q _18813_/Q vssd1 vssd1 vccd1 vccd1 _09126_/B sky130_fd_sc_hd__or3_4
XFILLER_31_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_175_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09054_ _09058_/A vssd1 vssd1 vccd1 vccd1 _09054_/Y sky130_fd_sc_hd__inv_2
XFILLER_135_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_1304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_173_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_172_1326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09956_ _12128_/A _09946_/X _09955_/X _09930_/X vssd1 vssd1 vccd1 vccd1 _09956_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_213_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09887_ _09902_/A _09887_/B vssd1 vssd1 vccd1 vccd1 _09979_/A sky130_fd_sc_hd__xnor2_4
XTAP_4127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10800_ _09160_/A _09160_/B _09165_/C _09170_/B _10770_/A _10812_/S vssd1 vssd1 vccd1
+ vccd1 _10800_/X sky130_fd_sc_hd__mux4_1
XTAP_2747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11780_ _11780_/A _11783_/A vssd1 vssd1 vccd1 vccd1 _11780_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_60_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10731_ _10731_/A _10731_/B vssd1 vssd1 vccd1 vccd1 _12100_/A sky130_fd_sc_hd__xnor2_2
XFILLER_214_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_213_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_194_wb_clk_i clkbuf_5_12_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18213_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_13450_ _13447_/A _13447_/B _13448_/Y _11720_/B _13449_/X vssd1 vssd1 vccd1 vccd1
+ _13450_/X sky130_fd_sc_hd__a221o_1
X_10662_ _10662_/A vssd1 vssd1 vccd1 vccd1 _10701_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_185_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_123_wb_clk_i clkbuf_5_25_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18434_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_16_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12401_ _18106_/Q _12401_/B vssd1 vssd1 vccd1 vccd1 _12403_/C sky130_fd_sc_hd__and2_1
XFILLER_22_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13381_ _17768_/A vssd1 vssd1 vccd1 vccd1 _13381_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_166_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10593_ _09720_/A _10589_/X _10592_/X _10582_/S vssd1 vssd1 vccd1 vccd1 _10593_/X
+ sky130_fd_sc_hd__a22o_1
X_15120_ _15266_/A _15134_/B vssd1 vssd1 vccd1 vccd1 _15132_/B sky130_fd_sc_hd__nor2_2
XFILLER_127_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12332_ _11415_/B _12330_/C _12347_/B vssd1 vssd1 vccd1 vccd1 _17883_/D sky130_fd_sc_hd__a21boi_1
XFILLER_5_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_181_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15051_ _15197_/A _15085_/B vssd1 vssd1 vccd1 vccd1 _15061_/B sky130_fd_sc_hd__nor2_1
XFILLER_147_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12263_ _12517_/A _12263_/B vssd1 vssd1 vccd1 vccd1 _12264_/A sky130_fd_sc_hd__and2_1
XFILLER_182_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14002_ _18925_/Q _13623_/A _13764_/A _18943_/Q vssd1 vssd1 vccd1 vccd1 _14002_/X
+ sky130_fd_sc_hd__a22o_1
X_11214_ _11214_/A vssd1 vssd1 vccd1 vccd1 _17815_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_141_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12194_ _17910_/Q _17909_/Q _17908_/Q _17907_/Q vssd1 vssd1 vccd1 vccd1 _12498_/A
+ sky130_fd_sc_hd__or4_2
X_18810_ _18811_/CLK _18810_/D vssd1 vssd1 vccd1 vccd1 _18810_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_6030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11145_ _17802_/Q vssd1 vssd1 vccd1 vccd1 _11922_/A sky130_fd_sc_hd__clkbuf_4
XTAP_6041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18741_ _18743_/CLK _18741_/D vssd1 vssd1 vccd1 vccd1 _18741_/Q sky130_fd_sc_hd__dfxtp_2
X_15953_ _16212_/A vssd1 vssd1 vccd1 vccd1 _16000_/A sky130_fd_sc_hd__clkbuf_2
XTAP_5340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11076_ _11590_/B vssd1 vssd1 vccd1 vccd1 _11368_/A sky130_fd_sc_hd__buf_2
XFILLER_209_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14904_ _15197_/A _14937_/B vssd1 vssd1 vccd1 vccd1 _14913_/B sky130_fd_sc_hd__nor2_1
X_10027_ _09136_/A _09126_/B _09131_/C _09136_/C _09986_/A _10025_/X vssd1 vssd1 vccd1
+ vccd1 _10027_/X sky130_fd_sc_hd__mux4_1
X_18672_ _18677_/CLK _18672_/D vssd1 vssd1 vccd1 vccd1 _18672_/Q sky130_fd_sc_hd__dfxtp_4
XTAP_5384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15884_ _18586_/Q _18550_/Q _15899_/S vssd1 vssd1 vccd1 vccd1 _15884_/X sky130_fd_sc_hd__mux2_1
XTAP_4650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17623_ _17687_/A _17663_/B vssd1 vssd1 vccd1 vccd1 _17623_/Y sky130_fd_sc_hd__nor2_2
XTAP_4683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14835_ _14872_/A _14838_/B vssd1 vssd1 vccd1 vccd1 _14835_/Y sky130_fd_sc_hd__nand2_1
XFILLER_5_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_224_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17554_ _14354_/X _16975_/X _17547_/X _17553_/X _14618_/X vssd1 vssd1 vccd1 vccd1
+ _18951_/D sky130_fd_sc_hd__o311a_1
X_14766_ _14948_/A vssd1 vssd1 vccd1 vccd1 _14814_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_63_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11978_ _11980_/A _11977_/Y _12015_/A vssd1 vssd1 vccd1 vccd1 _11978_/X sky130_fd_sc_hd__a21o_1
XFILLER_205_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_220_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16505_ _16510_/B _16502_/X _16504_/X _16496_/X vssd1 vssd1 vccd1 vccd1 _18696_/D
+ sky130_fd_sc_hd__o211a_1
X_10929_ _10927_/X _10928_/X _10935_/S vssd1 vssd1 vccd1 vccd1 _10929_/X sky130_fd_sc_hd__mux2_4
X_13717_ _18252_/Q _13716_/X _13654_/A _18243_/Q vssd1 vssd1 vccd1 vccd1 _13717_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_147_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14697_ _18265_/Q _14700_/B _14696_/Y _14692_/X vssd1 vssd1 vccd1 vccd1 _18265_/D
+ sky130_fd_sc_hd__o211a_1
X_17485_ _18970_/Q _18934_/Q _17495_/S vssd1 vssd1 vccd1 vccd1 _17485_/X sky130_fd_sc_hd__mux2_1
XFILLER_189_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19224_ _19224_/A _08932_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[24] sky130_fd_sc_hd__ebufn_8
X_16436_ _16447_/A _16439_/B vssd1 vssd1 vccd1 vccd1 _16436_/Y sky130_fd_sc_hd__nand2_1
XFILLER_32_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13648_ _13648_/A _13648_/B vssd1 vssd1 vccd1 vccd1 _13649_/C sky130_fd_sc_hd__nor2_1
XFILLER_32_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19155_ _19155_/A _08950_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[25] sky130_fd_sc_hd__ebufn_8
X_16367_ _16433_/A vssd1 vssd1 vccd1 vccd1 _16504_/C sky130_fd_sc_hd__clkbuf_2
X_13579_ _13579_/A vssd1 vssd1 vccd1 vccd1 _13580_/A sky130_fd_sc_hd__buf_8
XFILLER_121_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18106_ _18991_/CLK _18106_/D vssd1 vssd1 vccd1 vccd1 _18106_/Q sky130_fd_sc_hd__dfxtp_1
X_15318_ _15643_/A vssd1 vssd1 vccd1 vccd1 _15578_/A sky130_fd_sc_hd__clkbuf_2
X_16298_ _18681_/Q _18645_/Q _16304_/S vssd1 vssd1 vccd1 vccd1 _16298_/X sky130_fd_sc_hd__mux2_1
XFILLER_8_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19126__97 vssd1 vssd1 vccd1 vccd1 _19126__97/HI _19234_/A sky130_fd_sc_hd__conb_1
XFILLER_195_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_219_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18037_ _18094_/CLK _18037_/D vssd1 vssd1 vccd1 vccd1 _18037_/Q sky130_fd_sc_hd__dfxtp_1
X_15249_ _15253_/B _15246_/X _15248_/Y _15244_/X vssd1 vssd1 vccd1 vccd1 _18400_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_172_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_125_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09810_ _09810_/A _09810_/B _09810_/C vssd1 vssd1 vccd1 vccd1 _12106_/B sky130_fd_sc_hd__and3_1
XFILLER_99_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09741_ _18102_/Q _17981_/Q vssd1 vssd1 vccd1 vccd1 _09742_/B sky130_fd_sc_hd__xnor2_1
XFILLER_154_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_1204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18939_ _18939_/CLK _18939_/D vssd1 vssd1 vccd1 vccd1 _18939_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_189_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_1321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_227_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09672_ _09692_/A _09719_/B vssd1 vssd1 vccd1 vccd1 _10041_/A sky130_fd_sc_hd__xor2_4
XFILLER_27_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_223_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_223_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_270 _18396_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_1366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09106_ _18761_/Q _18760_/Q _18759_/Q vssd1 vssd1 vccd1 vccd1 _09109_/B sky130_fd_sc_hd__or3_4
XFILLER_175_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09037_ _09040_/A vssd1 vssd1 vccd1 vccd1 _09037_/Y sky130_fd_sc_hd__inv_2
XFILLER_184_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09939_ _09939_/A _09939_/B vssd1 vssd1 vccd1 vccd1 _10598_/A sky130_fd_sc_hd__xnor2_4
XFILLER_58_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12950_ _12961_/A vssd1 vssd1 vccd1 vccd1 _12950_/Y sky130_fd_sc_hd__inv_2
XFILLER_213_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11901_ _17791_/Q _17792_/Q vssd1 vssd1 vccd1 vccd1 _11927_/A sky130_fd_sc_hd__nor2_1
XTAP_3223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12881_ _17957_/Q _12881_/B vssd1 vssd1 vccd1 vccd1 _12886_/C sky130_fd_sc_hd__and2_1
XTAP_2500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11832_ _11905_/A _11832_/B _11832_/C vssd1 vssd1 vccd1 vccd1 _11859_/A sky130_fd_sc_hd__and3b_4
X_14620_ _14620_/A vssd1 vssd1 vccd1 vccd1 _17687_/A sky130_fd_sc_hd__buf_2
XTAP_3289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14551_ _16817_/A vssd1 vssd1 vccd1 vccd1 _15156_/A sky130_fd_sc_hd__buf_8
XTAP_1843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11763_ _11763_/A _11763_/B _11763_/C vssd1 vssd1 vccd1 vccd1 _11763_/X sky130_fd_sc_hd__and3_1
XTAP_1854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10714_ _10743_/A vssd1 vssd1 vccd1 vccd1 _10738_/A sky130_fd_sc_hd__buf_4
X_13502_ _13557_/B _13541_/B vssd1 vssd1 vccd1 vccd1 _13677_/A sky130_fd_sc_hd__nor2_1
XTAP_1887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14482_ _17420_/A vssd1 vssd1 vccd1 vccd1 _14491_/B sky130_fd_sc_hd__clkbuf_1
XTAP_1898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17270_ _17397_/B vssd1 vssd1 vccd1 vccd1 _17318_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_11694_ _17852_/Q _11704_/C _11339_/B _11703_/A vssd1 vssd1 vccd1 vccd1 _11694_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_105_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16221_ _16289_/A vssd1 vssd1 vccd1 vccd1 _16358_/C sky130_fd_sc_hd__buf_2
XFILLER_186_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13433_ _13649_/B _13649_/A _13648_/A _13635_/A vssd1 vssd1 vccd1 vccd1 _13436_/A
+ sky130_fd_sc_hd__and4b_1
X_10645_ _10661_/A _10661_/B vssd1 vssd1 vccd1 vccd1 _10770_/A sky130_fd_sc_hd__xnor2_4
XFILLER_9_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16152_ _18648_/Q _18612_/Q _16170_/S vssd1 vssd1 vccd1 vccd1 _16152_/X sky130_fd_sc_hd__mux2_1
XFILLER_127_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13364_ _17779_/Q _17780_/Q vssd1 vssd1 vccd1 vccd1 _17704_/B sky130_fd_sc_hd__and2b_1
XFILLER_158_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10576_ _09309_/D _10568_/X _10575_/X _10036_/A vssd1 vssd1 vccd1 vccd1 _10576_/X
+ sky130_fd_sc_hd__o211a_1
X_15103_ _15187_/A vssd1 vssd1 vccd1 vccd1 _15103_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_12315_ _12329_/A _11419_/X _11431_/B vssd1 vssd1 vccd1 vccd1 _12316_/C sky130_fd_sc_hd__o21a_1
X_16083_ _16082_/B _16080_/X _16082_/Y _16074_/X vssd1 vssd1 vccd1 vccd1 _18596_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_6_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_177_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13295_ _18054_/Q _18057_/Q _18056_/Q _18059_/Q vssd1 vssd1 vccd1 vccd1 _13297_/B
+ sky130_fd_sc_hd__or4_1
XFILLER_182_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15034_ _15058_/A _15038_/B vssd1 vssd1 vccd1 vccd1 _15034_/Y sky130_fd_sc_hd__nand2_1
X_12246_ _12246_/A _12269_/C vssd1 vssd1 vccd1 vccd1 _12246_/Y sky130_fd_sc_hd__nor2_1
XFILLER_29_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_91_wb_clk_i _18254_/CLK vssd1 vssd1 vccd1 vccd1 _18140_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_155_1321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_1354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12177_ _17847_/Q _12183_/B vssd1 vssd1 vccd1 vccd1 _12177_/X sky130_fd_sc_hd__and2_1
XFILLER_123_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_20_wb_clk_i clkbuf_5_4_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18899_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_96_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11128_ _13446_/A _11190_/A _11149_/S vssd1 vssd1 vccd1 vccd1 _11129_/A sky130_fd_sc_hd__mux2_1
XFILLER_111_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16985_ _14360_/X _16975_/X _16978_/X _16984_/Y _14618_/X vssd1 vssd1 vccd1 vccd1
+ _18809_/D sky130_fd_sc_hd__o311a_1
XFILLER_3_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18724_ _18724_/CLK _18724_/D vssd1 vssd1 vccd1 vccd1 _18724_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_27_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15936_ _15942_/B _15932_/X _15935_/X _15925_/X vssd1 vssd1 vccd1 vccd1 _18561_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_5170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11059_ _11059_/A vssd1 vssd1 vccd1 vccd1 _17786_/D sky130_fd_sc_hd__clkbuf_1
XTAP_5181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18655_ _18658_/CLK _18655_/D vssd1 vssd1 vccd1 vccd1 _18655_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_97_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15867_ _16019_/A _15892_/B vssd1 vssd1 vccd1 vccd1 _15876_/B sky130_fd_sc_hd__nor2_1
XTAP_4480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17606_ _17575_/X _17602_/Y _17603_/X _17605_/Y _18963_/Q vssd1 vssd1 vccd1 vccd1
+ _17607_/B sky130_fd_sc_hd__a32o_1
X_14818_ _14856_/A _15257_/B _14818_/C vssd1 vssd1 vccd1 vccd1 _14818_/X sky130_fd_sc_hd__or3_1
X_18586_ _18590_/CLK _18586_/D vssd1 vssd1 vccd1 vccd1 _18586_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_24_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15798_ _18564_/Q _18528_/Q _15809_/S vssd1 vssd1 vccd1 vccd1 _15798_/X sky130_fd_sc_hd__mux2_1
XFILLER_184_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_178_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17537_ _18984_/Q _18948_/Q _17543_/S vssd1 vssd1 vccd1 vccd1 _17537_/X sky130_fd_sc_hd__mux2_1
XFILLER_178_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14749_ _18313_/Q _18277_/Q _14756_/S vssd1 vssd1 vccd1 vccd1 _14749_/X sky130_fd_sc_hd__mux2_1
XFILLER_33_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_178_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_1347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17468_ _17468_/A vssd1 vssd1 vccd1 vccd1 _17512_/A sky130_fd_sc_hd__buf_2
XFILLER_220_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19207_ _19207_/A _08976_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[7] sky130_fd_sc_hd__ebufn_8
X_16419_ _16417_/B _16416_/X _16417_/Y _16418_/X vssd1 vssd1 vccd1 vccd1 _18674_/D
+ sky130_fd_sc_hd__o211a_1
X_17399_ _17437_/A _17538_/B _17399_/C vssd1 vssd1 vccd1 vccd1 _17399_/X sky130_fd_sc_hd__or3_1
XFILLER_160_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_1355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19138_ _19138_/A _09039_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[8] sky130_fd_sc_hd__ebufn_8
XFILLER_9_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_218_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_161_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_218_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09724_ _10070_/B vssd1 vssd1 vccd1 vccd1 _12063_/A sky130_fd_sc_hd__buf_2
XFILLER_210_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09655_ _10582_/S vssd1 vssd1 vccd1 vccd1 _12061_/A sky130_fd_sc_hd__buf_4
XFILLER_83_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_228_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_216_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09586_ _09586_/A _09586_/B vssd1 vssd1 vccd1 vccd1 _09587_/B sky130_fd_sc_hd__nand2_1
XFILLER_83_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_203_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_224_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_223_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_137_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_109_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10430_ _10561_/S vssd1 vssd1 vccd1 vccd1 _10430_/X sky130_fd_sc_hd__buf_4
XFILLER_137_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_183_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10361_ _09093_/A _09093_/B _09098_/C _09103_/B _09937_/X _12123_/A vssd1 vssd1 vccd1
+ vccd1 _10361_/X sky130_fd_sc_hd__mux4_2
XFILLER_164_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_178_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12100_ _12100_/A _12129_/A vssd1 vssd1 vccd1 vccd1 _12103_/B sky130_fd_sc_hd__xor2_1
XFILLER_124_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13080_ _13080_/A _17517_/A vssd1 vssd1 vccd1 vccd1 _13081_/A sky130_fd_sc_hd__and2_1
X_10292_ _09198_/A _09203_/B _10292_/S vssd1 vssd1 vccd1 vccd1 _10292_/X sky130_fd_sc_hd__mux2_1
XFILLER_128_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12031_ _12031_/A _13420_/A vssd1 vssd1 vccd1 vccd1 _12031_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_151_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_120_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16770_ _16769_/B _16767_/X _16769_/Y _16760_/X vssd1 vssd1 vccd1 vccd1 _18761_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_4_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13982_ _18358_/Q _13723_/X _13980_/X _13981_/X vssd1 vssd1 vccd1 vccd1 _13982_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_111_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_218_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15721_ _15719_/B _15718_/X _15719_/Y _15720_/X vssd1 vssd1 vccd1 vccd1 _18509_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_3020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_219_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12933_ _12933_/A _12933_/B vssd1 vssd1 vccd1 vccd1 _12933_/Y sky130_fd_sc_hd__nand2_1
XTAP_3031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_219_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_1355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18440_ _18443_/CLK _18440_/D vssd1 vssd1 vccd1 vccd1 _18440_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_18_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15652_ _15651_/B _15648_/X _15651_/Y _15640_/X vssd1 vssd1 vccd1 vccd1 _18491_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_18_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_222_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12864_ _12864_/A _12864_/B vssd1 vssd1 vccd1 vccd1 _17951_/D sky130_fd_sc_hd__nor2_1
XTAP_2341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_146_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14603_ _18243_/Q _14606_/B _14602_/X _14587_/X vssd1 vssd1 vccd1 vccd1 _18243_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_2363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18371_ _18374_/CLK _18371_/D vssd1 vssd1 vccd1 vccd1 _18371_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_15_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11815_ _17420_/A vssd1 vssd1 vccd1 vccd1 _17517_/A sky130_fd_sc_hd__clkbuf_4
XTAP_2374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15583_ _15633_/A _15583_/B vssd1 vssd1 vccd1 vccd1 _15583_/Y sky130_fd_sc_hd__nand2_1
XFILLER_15_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12795_ _17962_/Q vssd1 vssd1 vccd1 vccd1 _12795_/Y sky130_fd_sc_hd__inv_2
XTAP_2385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17322_ _17334_/A _17327_/B vssd1 vssd1 vccd1 vccd1 _17322_/Y sky130_fd_sc_hd__nand2_1
X_14534_ _18231_/Q _14545_/B _14532_/X _14533_/X vssd1 vssd1 vccd1 vccd1 _18231_/D
+ sky130_fd_sc_hd__o211a_1
X_11746_ _17915_/Q _17914_/Q vssd1 vssd1 vccd1 vccd1 _11761_/B sky130_fd_sc_hd__xnor2_2
XFILLER_30_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17253_ _17252_/B _17251_/X _17252_/Y _17241_/X vssd1 vssd1 vccd1 vccd1 _18875_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_41_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11677_ _11390_/X _11670_/X _11676_/X _11619_/X vssd1 vssd1 vccd1 vccd1 _11677_/X
+ sky130_fd_sc_hd__o22a_1
X_14465_ _14464_/A _14464_/B _12764_/X vssd1 vssd1 vccd1 vccd1 _14466_/B sky130_fd_sc_hd__o21ai_1
XFILLER_174_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16204_ _16959_/A vssd1 vssd1 vccd1 vccd1 _16794_/A sky130_fd_sc_hd__buf_4
X_13416_ _13416_/A vssd1 vssd1 vccd1 vccd1 _14355_/B sky130_fd_sc_hd__buf_2
X_10628_ _10640_/A _10656_/B vssd1 vssd1 vccd1 vccd1 _10661_/B sky130_fd_sc_hd__nor2_4
XFILLER_122_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14396_ _14396_/A vssd1 vssd1 vccd1 vccd1 _18190_/D sky130_fd_sc_hd__clkbuf_1
X_17184_ _17184_/A vssd1 vssd1 vccd1 vccd1 _17234_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_70_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16135_ _16734_/A _16150_/B vssd1 vssd1 vccd1 vccd1 _16147_/B sky130_fd_sc_hd__nor2_2
X_13347_ _13368_/A vssd1 vssd1 vccd1 vccd1 _13389_/B sky130_fd_sc_hd__buf_2
X_10559_ _09181_/C _09186_/B _10559_/S vssd1 vssd1 vccd1 vccd1 _10559_/X sky130_fd_sc_hd__mux2_1
XFILLER_128_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16066_ _16817_/A vssd1 vssd1 vccd1 vccd1 _16672_/A sky130_fd_sc_hd__buf_6
X_13278_ _13278_/A _13278_/B _13278_/C _13278_/D vssd1 vssd1 vccd1 vccd1 _13292_/A
+ sky130_fd_sc_hd__or4_1
XFILLER_29_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15017_ _15105_/A vssd1 vssd1 vccd1 vccd1 _15033_/S sky130_fd_sc_hd__clkbuf_2
X_12229_ _11606_/X _11614_/Y _12228_/Y _12233_/C _11614_/A vssd1 vssd1 vccd1 vccd1
+ _12230_/B sky130_fd_sc_hd__a32o_1
XFILLER_38_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_204_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_231_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16968_ _17032_/A _16972_/B vssd1 vssd1 vccd1 vccd1 _16968_/Y sky130_fd_sc_hd__nand2_1
XFILLER_83_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_226_wb_clk_i _17864_/CLK vssd1 vssd1 vccd1 vccd1 _17891_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_42_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18707_ _18710_/CLK _18707_/D vssd1 vssd1 vccd1 vccd1 _18707_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_225_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15919_ _16014_/A vssd1 vssd1 vccd1 vccd1 _15937_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_65_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16899_ _16903_/B _16895_/X _16898_/Y _16893_/X vssd1 vssd1 vccd1 vccd1 _18790_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_25_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09440_ _09440_/A vssd1 vssd1 vccd1 vccd1 _09440_/Y sky130_fd_sc_hd__inv_2
X_18638_ _18641_/CLK _18638_/D vssd1 vssd1 vccd1 vccd1 _18638_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_227_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_224_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_224_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09371_ _09371_/A _09371_/B _09371_/C vssd1 vssd1 vccd1 vccd1 _09427_/B sky130_fd_sc_hd__and3_2
X_18569_ _18571_/CLK _18569_/D vssd1 vssd1 vccd1 vccd1 _18569_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_206_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_220_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_212_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_162_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_1264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_221_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_192_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_158_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_3 _09034_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19110__81 vssd1 vssd1 vccd1 vccd1 _19110__81/HI _19218_/A sky130_fd_sc_hd__conb_1
XTAP_5928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_181_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09707_ _10102_/S vssd1 vssd1 vccd1 vccd1 _09708_/A sky130_fd_sc_hd__buf_2
XFILLER_114_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_228_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_215_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09638_ _09684_/A _09642_/B _09637_/X vssd1 vssd1 vccd1 vccd1 _09639_/B sky130_fd_sc_hd__o21a_1
XFILLER_83_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_203_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_128_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09569_ _10142_/A _09570_/B vssd1 vssd1 vccd1 vccd1 _09569_/X sky130_fd_sc_hd__and2_1
XFILLER_203_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_180_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11600_ _19034_/Q vssd1 vssd1 vccd1 vccd1 _11615_/A sky130_fd_sc_hd__inv_2
XFILLER_212_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_230_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12580_ _12580_/A vssd1 vssd1 vccd1 vccd1 _12582_/A sky130_fd_sc_hd__inv_2
XFILLER_196_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11531_ _11512_/C _11530_/X _19031_/Q vssd1 vssd1 vccd1 vccd1 _11531_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_8_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_212_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14250_ _18208_/Q vssd1 vssd1 vccd1 vccd1 _14464_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_11462_ _17886_/Q _11463_/B vssd1 vssd1 vccd1 vccd1 _12340_/A sky130_fd_sc_hd__or2_1
XFILLER_184_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13201_ _13201_/A vssd1 vssd1 vccd1 vccd1 _18056_/D sky130_fd_sc_hd__clkbuf_1
X_10413_ _10413_/A vssd1 vssd1 vccd1 vccd1 _10413_/X sky130_fd_sc_hd__buf_4
X_14181_ _18665_/Q _13539_/X _14175_/X _14180_/X vssd1 vssd1 vccd1 vccd1 _14181_/X
+ sky130_fd_sc_hd__a211o_1
X_11393_ _11655_/B _11539_/B _11790_/B vssd1 vssd1 vccd1 vccd1 _11393_/X sky130_fd_sc_hd__and3_1
XFILLER_137_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13132_ _13140_/A _18026_/Q vssd1 vssd1 vccd1 vccd1 _13133_/A sky130_fd_sc_hd__and2_1
X_10344_ _09136_/A _09126_/B _09131_/C _09136_/C _10307_/S _09905_/A vssd1 vssd1 vccd1
+ vccd1 _10345_/B sky130_fd_sc_hd__mux4_2
XFILLER_136_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_1321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17940_ _18151_/CLK _17940_/D vssd1 vssd1 vccd1 vccd1 _17940_/Q sky130_fd_sc_hd__dfxtp_2
X_13063_ _13063_/A _13063_/B vssd1 vssd1 vccd1 vccd1 _13063_/Y sky130_fd_sc_hd__nor2_1
XFILLER_97_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_215_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10275_ _09916_/X _10273_/X _09930_/A _10274_/X vssd1 vssd1 vccd1 vccd1 _10281_/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_152_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12014_ _11937_/C _12025_/A _12016_/B _11985_/D vssd1 vssd1 vccd1 vccd1 _12015_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_78_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17871_ _19030_/CLK _17871_/D vssd1 vssd1 vccd1 vccd1 _17871_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_79_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16822_ _18810_/Q _18774_/Q _16842_/S vssd1 vssd1 vccd1 vccd1 _16822_/X sky130_fd_sc_hd__mux2_1
XFILLER_78_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16753_ _16755_/B _16751_/X _16752_/Y _16740_/X vssd1 vssd1 vccd1 vccd1 _18757_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_93_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13965_ _18415_/Q _13642_/A _13764_/X _18439_/Q vssd1 vssd1 vccd1 vccd1 _13965_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_19_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15704_ _15751_/A _15708_/B vssd1 vssd1 vccd1 vccd1 _15704_/Y sky130_fd_sc_hd__nand2_1
XFILLER_206_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12916_ _12916_/A vssd1 vssd1 vccd1 vccd1 _17968_/D sky130_fd_sc_hd__clkbuf_1
X_16684_ _16686_/B _16680_/X _16681_/Y _16683_/X vssd1 vssd1 vccd1 vccd1 _18739_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_94_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13896_ _18598_/Q _13664_/X _13892_/X _13895_/X vssd1 vssd1 vccd1 vccd1 _13896_/X
+ sky130_fd_sc_hd__a211o_1
X_18423_ _18423_/CLK _18423_/D vssd1 vssd1 vccd1 vccd1 _18423_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_94_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15635_ _15677_/A vssd1 vssd1 vccd1 vccd1 _15696_/B sky130_fd_sc_hd__buf_2
XFILLER_61_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12847_ _12847_/A vssd1 vssd1 vccd1 vccd1 _12915_/B sky130_fd_sc_hd__clkbuf_2
XTAP_2171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_221_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18354_ _18356_/CLK _18354_/D vssd1 vssd1 vccd1 vccd1 _18354_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_72_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15566_ _15566_/A _15570_/B vssd1 vssd1 vccd1 vccd1 _15566_/Y sky130_fd_sc_hd__nand2_1
XFILLER_15_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12778_ _18004_/Q vssd1 vssd1 vccd1 vccd1 _13085_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_202_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17305_ _17303_/B _17302_/X _17303_/Y _17304_/X vssd1 vssd1 vccd1 vccd1 _18887_/D
+ sky130_fd_sc_hd__o211a_1
X_14517_ _14515_/Y _14516_/X _14436_/X vssd1 vssd1 vccd1 vccd1 _18229_/D sky130_fd_sc_hd__o21a_1
XFILLER_72_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18285_ _18317_/CLK _18285_/D vssd1 vssd1 vccd1 vccd1 _18285_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_30_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11729_ _11726_/Y _12509_/A _11729_/S vssd1 vssd1 vccd1 vccd1 _11729_/X sky130_fd_sc_hd__mux2_1
X_15497_ _15500_/B _15494_/X _15495_/Y _15496_/X vssd1 vssd1 vccd1 vccd1 _18454_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_174_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17236_ _18907_/Q _18871_/Q _17244_/S vssd1 vssd1 vccd1 vccd1 _17236_/X sky130_fd_sc_hd__mux2_1
X_14448_ _17564_/A _14448_/B vssd1 vssd1 vccd1 vccd1 _14449_/A sky130_fd_sc_hd__and2_1
XFILLER_156_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_190_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17167_ _18890_/Q _18854_/Q _17172_/S vssd1 vssd1 vccd1 vccd1 _17167_/X sky130_fd_sc_hd__mux2_1
XFILLER_31_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14379_ _18187_/Q _14375_/B _18188_/Q vssd1 vssd1 vccd1 vccd1 _14379_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_200_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16118_ _18640_/Q _18604_/Q _16145_/S vssd1 vssd1 vccd1 vccd1 _16118_/X sky130_fd_sc_hd__mux2_1
XFILLER_196_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17098_ _17098_/A vssd1 vssd1 vccd1 vccd1 _17114_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_116_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_118_1208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16049_ _16051_/B _16045_/X _16046_/Y _16048_/X vssd1 vssd1 vccd1 vccd1 _18589_/D
+ sky130_fd_sc_hd__o211a_1
X_08940_ _08941_/A vssd1 vssd1 vccd1 vccd1 _08940_/Y sky130_fd_sc_hd__inv_2
XFILLER_170_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_229_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_226_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_231_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_213_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09423_ _09427_/A _09423_/B vssd1 vssd1 vccd1 vccd1 _09450_/B sky130_fd_sc_hd__nand2_2
XFILLER_44_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_231_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_198_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09354_ _09354_/A _10389_/A _09354_/C _09354_/D vssd1 vssd1 vccd1 vccd1 _09355_/C
+ sky130_fd_sc_hd__and4_1
XFILLER_205_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_200_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09285_ _18863_/Q _18862_/Q _18861_/Q vssd1 vssd1 vccd1 vccd1 _09287_/C sky130_fd_sc_hd__or3_4
XFILLER_205_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_192_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19087__58 vssd1 vssd1 vccd1 vccd1 _19087__58/HI _19195_/A sky130_fd_sc_hd__conb_1
XFILLER_0_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_148_wb_clk_i clkbuf_5_26_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18275_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_5703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10060_ _10060_/A vssd1 vssd1 vccd1 vccd1 _10060_/X sky130_fd_sc_hd__clkbuf_4
XTAP_5714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_217_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13750_ _18783_/Q _13490_/A _13626_/A _18798_/Q vssd1 vssd1 vccd1 vccd1 _13750_/X
+ sky130_fd_sc_hd__a22o_1
X_10962_ _10962_/A _10962_/B vssd1 vssd1 vccd1 vccd1 _10962_/X sky130_fd_sc_hd__or2_1
XFILLER_18_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_216_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12701_ _12700_/Y _12707_/A _12699_/Y _12691_/B vssd1 vssd1 vccd1 vccd1 _12701_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_182_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13681_ _18534_/Q _13566_/A _13679_/X _13680_/X vssd1 vssd1 vccd1 vccd1 _13681_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_16_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10893_ _10891_/X _10892_/X _10893_/S vssd1 vssd1 vccd1 vccd1 _10893_/X sky130_fd_sc_hd__mux2_1
XFILLER_203_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_231_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15420_ _16019_/A _15448_/B vssd1 vssd1 vccd1 vccd1 _15431_/B sky130_fd_sc_hd__nor2_2
XFILLER_188_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12632_ _12632_/A _12632_/B vssd1 vssd1 vccd1 vccd1 _12632_/X sky130_fd_sc_hd__or2_1
XFILLER_203_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_231_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_223_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15351_ _18458_/Q _18422_/Q _15356_/S vssd1 vssd1 vccd1 vccd1 _15351_/X sky130_fd_sc_hd__mux2_1
XFILLER_212_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12563_ _12594_/B _17920_/Q vssd1 vssd1 vccd1 vccd1 _12563_/Y sky130_fd_sc_hd__nand2_1
XFILLER_15_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_223_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11514_ _17870_/Q vssd1 vssd1 vccd1 vccd1 _12279_/A sky130_fd_sc_hd__clkbuf_2
X_14302_ _15463_/B vssd1 vssd1 vccd1 vccd1 _15145_/A sky130_fd_sc_hd__buf_4
X_18070_ _18072_/CLK _18070_/D vssd1 vssd1 vccd1 vccd1 _18070_/Q sky130_fd_sc_hd__dfxtp_1
X_15282_ _15301_/A _15286_/B vssd1 vssd1 vccd1 vccd1 _15282_/Y sky130_fd_sc_hd__nand2_1
X_12494_ _12495_/A _12495_/B _12495_/C _12495_/D vssd1 vssd1 vccd1 vccd1 _12496_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_7_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17021_ _17023_/B _17017_/X _17018_/Y _17020_/X vssd1 vssd1 vccd1 vccd1 _18817_/D
+ sky130_fd_sc_hd__o211a_1
X_11445_ _11661_/A _11396_/B _11413_/Y _11436_/Y _11444_/X vssd1 vssd1 vccd1 vccd1
+ _11445_/X sky130_fd_sc_hd__a41o_1
X_14233_ _14233_/A _18206_/Q vssd1 vssd1 vccd1 vccd1 _14463_/B sky130_fd_sc_hd__nand2_1
XFILLER_171_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14164_ _18983_/Q _13617_/X _14162_/X _14163_/X vssd1 vssd1 vccd1 vccd1 _14164_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_153_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11376_ _11376_/A _11376_/B vssd1 vssd1 vccd1 vccd1 _11377_/A sky130_fd_sc_hd__nand2_1
XFILLER_166_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_217_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13115_ _13115_/A vssd1 vssd1 vccd1 vccd1 _18017_/D sky130_fd_sc_hd__clkbuf_1
X_10327_ _10338_/A _10323_/X _10326_/X _09921_/X vssd1 vssd1 vccd1 vccd1 _10327_/X
+ sky130_fd_sc_hd__a22o_1
X_14095_ _18446_/Q _14015_/A _13515_/X _18422_/Q _14094_/X vssd1 vssd1 vccd1 vccd1
+ _14095_/X sky130_fd_sc_hd__a221o_2
XFILLER_152_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18972_ _18972_/CLK _18972_/D vssd1 vssd1 vccd1 vccd1 _18972_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13046_ _13049_/A _13046_/B vssd1 vssd1 vccd1 vccd1 _13047_/A sky130_fd_sc_hd__and2_1
X_17923_ _17926_/CLK _17923_/D vssd1 vssd1 vccd1 vccd1 _17923_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_79_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10258_ _10191_/A _10258_/B vssd1 vssd1 vccd1 vccd1 _10258_/X sky130_fd_sc_hd__and2b_1
XFILLER_112_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_230_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17854_ _17895_/CLK _17854_/D vssd1 vssd1 vccd1 vccd1 _17854_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_113_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_1176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10189_ _18120_/Q _10189_/B vssd1 vssd1 vccd1 vccd1 _10191_/A sky130_fd_sc_hd__xnor2_1
X_16805_ _17410_/A _16976_/B vssd1 vssd1 vccd1 vccd1 _16879_/A sky130_fd_sc_hd__or2_1
XFILLER_82_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17785_ _17817_/CLK _17785_/D vssd1 vssd1 vccd1 vccd1 _17785_/Q sky130_fd_sc_hd__dfxtp_1
X_14997_ _15145_/C _15145_/A _15145_/B vssd1 vssd1 vccd1 vccd1 _15064_/A sky130_fd_sc_hd__or3b_4
XFILLER_93_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16736_ _16736_/A _16736_/B _16773_/C vssd1 vssd1 vccd1 vccd1 _16736_/X sky130_fd_sc_hd__or3_1
X_13948_ _18499_/Q _13579_/A _13624_/A _18493_/Q vssd1 vssd1 vccd1 vccd1 _13948_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_75_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_223_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_222_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_207_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16667_ _18735_/Q _16670_/B _16666_/X _16659_/X vssd1 vssd1 vccd1 vccd1 _18735_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_61_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13879_ _18883_/Q _13869_/A _13861_/A _18907_/Q _13878_/X vssd1 vssd1 vccd1 vccd1
+ _13879_/X sky130_fd_sc_hd__a221o_1
XFILLER_62_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18406_ _18406_/CLK _18406_/D vssd1 vssd1 vccd1 vccd1 _18406_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_61_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15618_ _15633_/A _15618_/B vssd1 vssd1 vccd1 vccd1 _15618_/Y sky130_fd_sc_hd__nand2_1
XFILLER_179_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16598_ _18755_/Q _18719_/Q _16598_/S vssd1 vssd1 vccd1 vccd1 _16598_/X sky130_fd_sc_hd__mux2_1
XFILLER_50_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18337_ _18373_/CLK _18337_/D vssd1 vssd1 vccd1 vccd1 _18337_/Q sky130_fd_sc_hd__dfxtp_1
X_15549_ _15568_/A vssd1 vssd1 vccd1 vccd1 _15565_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_187_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09070_ _09070_/A vssd1 vssd1 vccd1 vccd1 _19178_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_136_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18268_ _18275_/CLK _18268_/D vssd1 vssd1 vccd1 vccd1 _18268_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_129_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17219_ _17304_/A vssd1 vssd1 vccd1 vccd1 _17219_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_190_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18199_ _18203_/CLK _18199_/D vssd1 vssd1 vccd1 vccd1 _18199_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_190_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_226_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09972_ _09972_/A _09972_/B vssd1 vssd1 vccd1 vccd1 _09972_/X sky130_fd_sc_hd__or2_1
XFILLER_226_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_218_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_217_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_225_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09406_ _18308_/Q _18307_/Q _18306_/Q vssd1 vssd1 vccd1 vccd1 _09408_/C sky130_fd_sc_hd__or3_2
XFILLER_80_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09337_ _09337_/A _09337_/B _09337_/C _09337_/D vssd1 vssd1 vccd1 vccd1 _09338_/C
+ sky130_fd_sc_hd__and4_1
XFILLER_200_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09268_ _18968_/Q _18967_/Q _18966_/Q vssd1 vssd1 vccd1 vccd1 _09270_/C sky130_fd_sc_hd__or3_2
XFILLER_103_1318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_181_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09199_ _18566_/Q _18565_/Q _18564_/Q vssd1 vssd1 vccd1 vccd1 _09203_/A sky130_fd_sc_hd__or3_2
XFILLER_147_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11230_ _11232_/A _11232_/C _11221_/X vssd1 vssd1 vccd1 vccd1 _11231_/B sky130_fd_sc_hd__o21ai_1
XFILLER_107_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_175_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11161_ _17818_/Q _17819_/Q _17821_/Q _17820_/Q vssd1 vssd1 vccd1 vccd1 _11164_/C
+ sky130_fd_sc_hd__or4b_2
XFILLER_84_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10112_ _18118_/Q _10114_/B vssd1 vssd1 vccd1 vccd1 _10120_/A sky130_fd_sc_hd__nand2_1
XFILLER_161_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11092_ _11092_/A vssd1 vssd1 vccd1 vccd1 _17792_/D sky130_fd_sc_hd__clkbuf_1
XTAP_5511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_216_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14920_ _18318_/Q _14924_/B _14919_/X _14902_/X vssd1 vssd1 vccd1 vccd1 _18318_/D
+ sky130_fd_sc_hd__o211a_1
X_10043_ _09219_/A _09209_/C _10795_/A _09214_/C _10004_/B _10025_/X vssd1 vssd1 vccd1
+ vccd1 _10044_/B sky130_fd_sc_hd__mux4_1
XTAP_5544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_212_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14851_ _15145_/B _15145_/C _15145_/A vssd1 vssd1 vccd1 vccd1 _14918_/A sky130_fd_sc_hd__or3b_4
XTAP_5599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13802_ _18357_/Q _13742_/X _13800_/X _13801_/X vssd1 vssd1 vccd1 vccd1 _13802_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_35_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17570_ _17570_/A vssd1 vssd1 vccd1 vccd1 _18955_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14782_ _14793_/A _15220_/B _14818_/C vssd1 vssd1 vccd1 vccd1 _14782_/X sky130_fd_sc_hd__or3_1
XFILLER_28_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11994_ _11541_/B _11499_/C _11922_/B vssd1 vssd1 vccd1 vccd1 _13518_/B sky130_fd_sc_hd__a21o_4
XFILLER_44_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16521_ _16521_/A vssd1 vssd1 vccd1 vccd1 _16572_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_186_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13733_ _13733_/A vssd1 vssd1 vccd1 vccd1 _13733_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_205_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_189_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10945_ _10941_/X _10943_/X _10944_/X _10010_/X _09709_/X vssd1 vssd1 vccd1 vccd1
+ _10945_/X sky130_fd_sc_hd__a221o_1
XFILLER_182_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_45_wb_clk_i clkbuf_5_18_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18811_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_95_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16452_ _16745_/A _16452_/B vssd1 vssd1 vccd1 vccd1 _16464_/B sky130_fd_sc_hd__nor2_2
XFILLER_231_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13664_ _13664_/A vssd1 vssd1 vccd1 vccd1 _13664_/X sky130_fd_sc_hd__buf_4
XFILLER_16_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10876_ _09402_/A _09392_/B _10882_/S vssd1 vssd1 vccd1 vccd1 _10876_/X sky130_fd_sc_hd__mux2_1
XFILLER_147_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15403_ _15445_/A _15403_/B vssd1 vssd1 vccd1 vccd1 _15403_/Y sky130_fd_sc_hd__nand2_1
XPHY_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12615_ _17929_/Q _17926_/Q vssd1 vssd1 vccd1 vccd1 _12616_/A sky130_fd_sc_hd__xnor2_1
X_19171_ _19171_/A _09019_/Y vssd1 vssd1 vccd1 vccd1 io_out[9] sky130_fd_sc_hd__ebufn_8
XFILLER_223_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16383_ _16473_/A vssd1 vssd1 vccd1 vccd1 _16400_/S sky130_fd_sc_hd__buf_2
XPHY_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13595_ _13705_/A vssd1 vssd1 vccd1 vccd1 _13596_/A sky130_fd_sc_hd__buf_6
XPHY_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18122_ _18130_/CLK _18122_/D vssd1 vssd1 vccd1 vccd1 _18122_/Q sky130_fd_sc_hd__dfxtp_2
X_15334_ _18454_/Q _18418_/Q _15334_/S vssd1 vssd1 vccd1 vccd1 _15334_/X sky130_fd_sc_hd__mux2_1
XPHY_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_223_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12546_ _12635_/A vssd1 vssd1 vccd1 vccd1 _12569_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_8_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_185_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18053_ _18068_/CLK _18053_/D vssd1 vssd1 vccd1 vccd1 _18053_/Q sky130_fd_sc_hd__dfxtp_1
X_15265_ _15263_/B _15262_/X _15263_/Y _15264_/X vssd1 vssd1 vccd1 vccd1 _18404_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_145_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12477_ _12477_/A _12477_/B _12477_/C _12477_/D vssd1 vssd1 vccd1 vccd1 _12499_/D
+ sky130_fd_sc_hd__nor4_2
XFILLER_126_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17004_ _17010_/B _17002_/X _17003_/X _16999_/X vssd1 vssd1 vccd1 vccd1 _18813_/D
+ sky130_fd_sc_hd__o211a_1
X_14216_ _14216_/A _14216_/B vssd1 vssd1 vccd1 vccd1 _14342_/A sky130_fd_sc_hd__nor2_1
X_11428_ _17883_/Q _11428_/B vssd1 vssd1 vccd1 vccd1 _11428_/Y sky130_fd_sc_hd__nand2_1
X_15196_ _15195_/B _15193_/X _15195_/Y _15187_/X vssd1 vssd1 vccd1 vccd1 _18386_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_6_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_158_1363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14147_ _18575_/Q _13523_/A _13598_/X _18557_/Q vssd1 vssd1 vccd1 vccd1 _14147_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_154_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11359_ _17796_/Q _11359_/B vssd1 vssd1 vccd1 vccd1 _11506_/B sky130_fd_sc_hd__and2_1
XFILLER_125_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_98_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14078_ _18731_/Q _13838_/A _14076_/X _14077_/X vssd1 vssd1 vccd1 vccd1 _14078_/X
+ sky130_fd_sc_hd__a211o_1
X_18955_ _18959_/CLK _18955_/D vssd1 vssd1 vccd1 vccd1 _18955_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_140_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17906_ _17907_/CLK _17906_/D vssd1 vssd1 vccd1 vccd1 _17906_/Q sky130_fd_sc_hd__dfxtp_1
X_13029_ _12982_/A _13025_/X _13028_/X _13011_/X vssd1 vssd1 vccd1 vccd1 _17987_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_117_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18886_ _18899_/CLK _18886_/D vssd1 vssd1 vccd1 vccd1 _18886_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_6_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17837_ _18992_/CLK _17837_/D vssd1 vssd1 vccd1 vccd1 _17837_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_55_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_227_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17768_ _17768_/A _17768_/B _17768_/C vssd1 vssd1 vccd1 vccd1 _17769_/A sky130_fd_sc_hd__and3_1
XFILLER_214_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_1304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16719_ _18784_/Q _18748_/Q _16742_/S vssd1 vssd1 vccd1 vccd1 _16719_/X sky130_fd_sc_hd__mux2_1
XFILLER_19_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17699_ _18987_/Q _17698_/Y _17705_/S vssd1 vssd1 vccd1 vccd1 _17700_/A sky130_fd_sc_hd__mux2_1
XFILLER_179_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_222_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_206_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09122_ _18839_/Q _18838_/Q _18837_/Q vssd1 vssd1 vccd1 vccd1 _09126_/A sky130_fd_sc_hd__or3_4
XFILLER_148_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_202_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09053_ _09053_/A vssd1 vssd1 vccd1 vccd1 _09058_/A sky130_fd_sc_hd__buf_12
XFILLER_175_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19057__28 vssd1 vssd1 vccd1 vccd1 _19057__28/HI _19151_/A sky130_fd_sc_hd__conb_1
XFILLER_131_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09955_ _14240_/B _09949_/X _09954_/X _10305_/S vssd1 vssd1 vccd1 vccd1 _09955_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_132_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_213_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09886_ _09974_/A vssd1 vssd1 vccd1 vccd1 _10370_/S sky130_fd_sc_hd__clkbuf_4
XTAP_870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_213_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_198_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_198_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10730_ _10664_/A _10727_/X _10729_/X _10818_/A vssd1 vssd1 vccd1 vccd1 _10730_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_199_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_213_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_185_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10661_ _10661_/A _10661_/B vssd1 vssd1 vccd1 vccd1 _10662_/A sky130_fd_sc_hd__xor2_4
XFILLER_213_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_201_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12400_ _18106_/Q _12401_/B vssd1 vssd1 vccd1 vccd1 _12409_/B sky130_fd_sc_hd__nor2_1
XFILLER_220_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13380_ _13380_/A vssd1 vssd1 vccd1 vccd1 _18112_/D sky130_fd_sc_hd__clkbuf_1
X_10592_ _10590_/X _10591_/X _10893_/S vssd1 vssd1 vccd1 vccd1 _10592_/X sky130_fd_sc_hd__mux2_1
XFILLER_222_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_1178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12331_ _12331_/A vssd1 vssd1 vccd1 vccd1 _17882_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_108_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_163_wb_clk_i clkbuf_5_11_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18068_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_5_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15050_ _15049_/B _15048_/X _15049_/Y _15046_/X vssd1 vssd1 vccd1 vccd1 _18350_/D
+ sky130_fd_sc_hd__o211a_1
X_12262_ _12261_/Y _12261_/A _12270_/A vssd1 vssd1 vccd1 vccd1 _12263_/B sky130_fd_sc_hd__mux2_1
X_11213_ _11215_/B _11243_/A vssd1 vssd1 vccd1 vccd1 _11214_/A sky130_fd_sc_hd__and2b_1
X_14001_ _18931_/Q _13666_/X _13781_/X _18928_/Q _14000_/X vssd1 vssd1 vccd1 vccd1
+ _14001_/X sky130_fd_sc_hd__a221o_1
XFILLER_135_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12193_ _17893_/Q _17892_/Q _12352_/B _12193_/D vssd1 vssd1 vccd1 vccd1 _12198_/A
+ sky130_fd_sc_hd__or4_1
XFILLER_150_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11144_ _11144_/A vssd1 vssd1 vccd1 vccd1 _17801_/D sky130_fd_sc_hd__clkbuf_1
XTAP_6020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18740_ _18743_/CLK _18740_/D vssd1 vssd1 vccd1 vccd1 _18740_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_95_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15952_ _17222_/A vssd1 vssd1 vccd1 vccd1 _16212_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_153_1260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11075_ _11975_/A vssd1 vssd1 vccd1 vccd1 _11590_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_110_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14903_ _14900_/B _14899_/X _14900_/Y _14902_/X vssd1 vssd1 vccd1 vccd1 _18314_/D
+ sky130_fd_sc_hd__o211a_1
X_10026_ _09126_/A _09136_/B _09131_/A _09126_/D _10956_/B _10025_/X vssd1 vssd1 vccd1
+ vccd1 _10026_/X sky130_fd_sc_hd__mux4_1
XFILLER_49_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18671_ _18677_/CLK _18671_/D vssd1 vssd1 vccd1 vccd1 _18671_/Q sky130_fd_sc_hd__dfxtp_4
XTAP_5374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15883_ _15883_/A vssd1 vssd1 vccd1 vccd1 _15899_/S sky130_fd_sc_hd__clkbuf_2
XTAP_4640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17622_ _14360_/X _14612_/A _17547_/A _17621_/X _17556_/X vssd1 vssd1 vccd1 vccd1
+ _18968_/D sky130_fd_sc_hd__o311a_1
XFILLER_224_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19071__42 vssd1 vssd1 vccd1 vccd1 _19071__42/HI _19165_/A sky130_fd_sc_hd__conb_1
XTAP_4673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14834_ _18334_/Q _18298_/Q _14848_/S vssd1 vssd1 vccd1 vccd1 _14834_/X sky130_fd_sc_hd__mux2_1
XTAP_4684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17553_ _17548_/Y _17552_/X _18951_/Q vssd1 vssd1 vccd1 vccd1 _17553_/X sky130_fd_sc_hd__a21o_1
XTAP_3983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14765_ _18317_/Q _18281_/Q _14787_/S vssd1 vssd1 vccd1 vccd1 _14765_/X sky130_fd_sc_hd__mux2_1
XTAP_3994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11977_ _11985_/A _12025_/D vssd1 vssd1 vccd1 vccd1 _11977_/Y sky130_fd_sc_hd__nor2_1
XFILLER_32_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16504_ _16555_/A _16796_/B _16504_/C vssd1 vssd1 vccd1 vccd1 _16504_/X sky130_fd_sc_hd__or3_1
XFILLER_72_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13716_ _13760_/A vssd1 vssd1 vccd1 vccd1 _13716_/X sky130_fd_sc_hd__buf_4
XFILLER_17_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_204_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10928_ _09332_/A _09327_/A _09337_/B _10782_/A _10462_/X _10450_/S vssd1 vssd1 vccd1
+ vccd1 _10928_/X sky130_fd_sc_hd__mux4_1
X_17484_ _17489_/B _17482_/X _17483_/X _17478_/X vssd1 vssd1 vccd1 vccd1 _18933_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_220_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14696_ _14750_/A _14700_/B vssd1 vssd1 vccd1 vccd1 _14696_/Y sky130_fd_sc_hd__nand2_1
XFILLER_16_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19223_ _19223_/A _08957_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[23] sky130_fd_sc_hd__ebufn_8
X_16435_ _18678_/Q _16439_/B _16434_/X _16418_/X vssd1 vssd1 vccd1 vccd1 _18678_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_20_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_177_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13647_ _18912_/Q _13575_/A _13576_/A _18903_/Q _13646_/X vssd1 vssd1 vccd1 vccd1
+ _13647_/X sky130_fd_sc_hd__a221o_1
XFILLER_220_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10859_ _10857_/X _10858_/X _10859_/S vssd1 vssd1 vccd1 vccd1 _10859_/X sky130_fd_sc_hd__mux2_1
XFILLER_13_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19154_ _19154_/A _08948_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[24] sky130_fd_sc_hd__ebufn_8
XPHY_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16366_ _17549_/A _16366_/B vssd1 vssd1 vccd1 vccd1 _16433_/A sky130_fd_sc_hd__or2_1
XFILLER_9_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13578_ _13772_/A vssd1 vssd1 vccd1 vccd1 _13579_/A sky130_fd_sc_hd__buf_6
XFILLER_121_1215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18105_ _18988_/CLK _18105_/D vssd1 vssd1 vccd1 vccd1 _18105_/Q sky130_fd_sc_hd__dfxtp_1
X_15317_ _18451_/Q _18415_/Q _15334_/S vssd1 vssd1 vccd1 vccd1 _15317_/X sky130_fd_sc_hd__mux2_1
XFILLER_121_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12529_ _12591_/A vssd1 vssd1 vccd1 vccd1 _12529_/X sky130_fd_sc_hd__clkbuf_2
X_16297_ _16734_/A _16307_/B vssd1 vssd1 vccd1 vccd1 _16305_/B sky130_fd_sc_hd__nor2_1
XFILLER_173_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_1319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18036_ _18094_/CLK _18036_/D vssd1 vssd1 vccd1 vccd1 _18036_/Q sky130_fd_sc_hd__dfxtp_1
X_15248_ _15301_/A _15253_/B vssd1 vssd1 vccd1 vccd1 _15248_/Y sky130_fd_sc_hd__nand2_1
XFILLER_114_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15179_ _15182_/B _15177_/X _15178_/Y _15166_/X vssd1 vssd1 vccd1 vccd1 _18382_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_125_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_132_1300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09740_ _09752_/A _09752_/B vssd1 vssd1 vccd1 vccd1 _09753_/A sky130_fd_sc_hd__nand2_1
XFILLER_228_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18938_ _18965_/CLK _18938_/D vssd1 vssd1 vccd1 vccd1 _18938_/Q sky130_fd_sc_hd__dfxtp_2
.ends

